# 5 3.10862e-13
(0,127) x (0,63)
[ (-1.1279e-24,2.01968e-24) (4.19397e-23,1.79351e-23) (1.73698e-22,-3.41121e-22) (-6.33818e-21,-2.23519e-21) (-2.38881e-20,5.01933e-20) (8.19163e-19,2.38788e-19) (2.94809e-18,-6.40686e-18) (-8.91874e-17,-2.19115e-17) (-3.26708e-16,7.0215e-16) (8.05201e-15,1.77313e-15) (3.19242e-14,-6.50326e-14) (-5.92704e-13,-1.33281e-13) (-2.66417e-12,4.97977e-12) (3.49173e-11,9.62908e-12) (1.82996e-10,-3.06149e-10) (-1.61109e-09,-6.4105e-10) (-9.97261e-09,1.45341e-08) (5.65156e-08,3.55994e-08) (4.15986e-07,-5.0558e-07) (-1.42706e-06,-1.49077e-06) (-1.27157e-05,1.19581e-05) (2.29398e-05,4.28579e-05) (0.000264874,-0.000170073) (-0.000166072,-0.00074997) (-0.00328464,0.00109743) (-0.000303464,0.00644028) (0.019973,-4.05013e-05) (0.00829977,-0.0140226) (-0.041913,-0.0222868) (-0.033392,-0.0526095) (-0.0232642,0.024182) (-0.11808,-0.0773275) (0.0495418,-0.0929664) (-0.0764215,0.0218445) (-0.103991,-0.15112) (-0.0409774,-0.0402693) (-0.139562,0.00488763) (0.1307,-0.00589284) (0.0381049,-0.00942995) (-0.0545768,0.0383814) (0.00913011,-0.0244498) (0.00295171,0.000611823) (-0.00125472,0.00689356) (0.000257942,-0.0018131) (-0.000179453,-0.000666168) (-3.82061e-05,0.000186583) (1.32336e-05,3.70022e-05) (4.87958e-06,-8.92209e-06) (-4.8295e-07,-1.23003e-06) (-2.85976e-07,2.5311e-07) (1.46232e-08,2.74351e-08) (1.00704e-08,-5.06837e-09) (-5.88222e-10,-3.47082e-10) (-2.40554e-10,8.79659e-11) (1.97787e-11,-3.00167e-12) (4.15327e-12,-1.34412e-12) (-4.92295e-13,1.98382e-13) (-5.80376e-14,3.61942e-14) (1.17467e-14,-8.25285e-15) (8.83068e-16,-2.24504e-16) (-3.24775e-16,2.41945e-16) (-1.41453e-17,-1.99798e-17) (7.45674e-18,-4.53434e-18) (1.85135e-19,6.74364e-19) 
  (-2.58628e-25,4.69045e-24) (7.22413e-23,-1.20408e-23) (-2.33771e-24,-7.577e-22) (-1.04439e-20,2.29564e-21) (5.61604e-21,1.06672e-19) (1.30214e-18,-3.37903e-19) (-1.20107e-18,-1.30259e-17) (-1.38268e-16,3.86569e-17) (1.60809e-16,1.36959e-15) (1.23563e-14,-3.36296e-15) (-1.53045e-14,-1.22435e-13) (-9.18571e-13,2.09447e-13) (1.03404e-12,9.13335e-12) (5.60922e-11,-7.7828e-12) (-4.48058e-11,-5.54157e-10) (-2.76825e-09,7.46514e-13) (6.60445e-10,2.64412e-08) (1.07693e-07,1.99949e-08) (5.91543e-08,-9.50474e-07) (-3.16182e-06,-1.31973e-06) (-4.7512e-06,2.43458e-05) (6.48081e-05,4.60093e-05) (0.000161418,-0.00041) (-0.000804641,-0.000907126) (-0.0027358,0.00395238) (0.00451322,0.00870428) (0.0208185,-0.0174494) (0.00260426,-0.0259555) (-0.0559995,0.0164893) (-0.0955054,-0.0255016) (0.00772521,0.0318448) (-0.188366,0.0607176) (-0.0633008,-0.151498) (-0.0284857,0.0931577) (-0.254836,-0.0315074) (-0.0824081,-0.00393345) (-0.166569,0.155227) (0.111949,-0.120567) (0.0479545,-0.0668111) (-0.0195827,0.0925825) (-0.0149218,-0.0275105) (0.00306002,-0.00462903) (0.00553533,0.00801969) (-0.00120157,-0.00169806) (-0.000924995,-0.000550904) (0.000107622,0.000213491) (5.89121e-05,2.98751e-05) (-1.76601e-06,-1.35978e-05) (-2.08793e-06,-1.16109e-06) (-1.07261e-07,5.37629e-07) (5.07051e-08,3.0999e-08) (6.67421e-09,-1.52928e-08) (-1.05406e-09,-3.08244e-10) (-1.78899e-10,3.46343e-10) (1.80453e-11,-1.07505e-11) (2.95863e-12,-6.27066e-12) (-3.06918e-13,4.94082e-13) (-1.94564e-14,1.14397e-13) (4.30839e-15,-1.72998e-14) (4.64585e-16,-1.58514e-15) (-8.64353e-17,5.31076e-16) (-2.80478e-17,6.54305e-18) (2.24609e-18,-1.15889e-17) (7.51711e-19,2.24693e-19) 
  (2.93972e-24,5.65652e-24) (6.55149e-23,-5.31184e-23) (-5.17279e-22,-8.60591e-22) (-9.14818e-21,8.13872e-21) (7.72571e-20,1.13973e-19) (1.11509e-18,-1.0537e-18) (-9.76628e-18,-1.30655e-17) (-1.18041e-16,1.13249e-16) (1.03579e-15,1.29084e-15) (1.07869e-14,-9.90731e-15) (-9.09497e-14,-1.09119e-13) (-8.4308e-13,6.8872e-13) (6.49074e-12,7.79652e-12) (5.54494e-11,-3.68253e-11) (-3.66717e-10,-4.61786e-10) (-2.99018e-09,1.43849e-09) (1.57662e-08,2.20415e-08) (1.27489e-07,-3.6851e-08) (-4.84675e-07,-8.16319e-07) (-4.09562e-06,4.04601e-07) (9.59065e-06,2.22878e-05) (9.25793e-05,8.56068e-06) (-9.78222e-05,-0.00041493) (-0.00131244,-0.000395024) (0.000121364,0.00461046) (0.00933009,0.00541652) (0.00456374,-0.0249053) (-0.0131521,-0.0276594) (-0.0224287,0.0421348) (-0.0947736,0.0522682) (0.0180259,0.000588464) (-0.0698052,0.181756) (-0.17235,-0.0514526) (0.0569581,0.0630104) (-0.190347,0.165704) (-0.0605134,0.0514156) (-0.0221811,0.255728) (-0.0068287,-0.138408) (-0.011948,-0.106832) (0.0484894,0.0785714) (-0.0256871,-0.00439438) (-0.00272035,-0.00649451) (0.009297,0.00164442) (-0.00154976,-0.000327556) (-0.00111972,0.000271425) (0.000186653,9.69673e-05) (7.1939e-05,-2.11149e-05) (-8.76756e-06,-1.004e-05) (-2.80976e-06,5.49235e-07) (2.31416e-07,5.15758e-07) (7.56048e-08,-4.56019e-09) (-4.30082e-09,-1.6942e-08) (-1.4176e-09,1.63047e-10) (9.30476e-11,4.01838e-10) (1.47208e-11,-1.17122e-11) (-2.39065e-12,-7.12415e-12) (-3.39873e-14,4.25266e-13) (7.69977e-14,1.06136e-13) (-6.17351e-15,-1.38657e-14) (-1.18559e-15,-1.65232e-15) (2.73989e-16,4.16025e-16) (-3.14041e-18,2.88489e-17) (-6.48612e-18,-9.1083e-18) (4.3536e-19,-4.67863e-19) 
  (5.7751e-24,3.43126e-24) (3.1634e-23,-7.5248e-23) (-9.23296e-22,-4.75344e-22) (-4.04105e-21,1.10467e-20) (1.27041e-19,5.71062e-20) (4.59665e-19,-1.39151e-18) (-1.49257e-17,-5.92664e-18) (-4.76374e-17,1.4846e-16) (1.48421e-15,5.32819e-16) (4.55778e-15,-1.32302e-14) (-1.23538e-13,-4.17339e-14) (-3.96313e-13,9.6962e-13) (8.48287e-12,2.85656e-12) (2.99142e-11,-5.73466e-11) (-4.70945e-10,-1.69523e-10) (-1.85018e-09,2.6696e-09) (2.05291e-08,8.51436e-09) (8.88325e-08,-9.44391e-08) (-6.73697e-07,-3.47088e-07) (-3.14889e-06,2.40761e-06) (1.57025e-05,1.07565e-05) (7.75555e-05,-4.04753e-05) (-0.000239704,-0.000228577) (-0.00120026,0.000370954) (0.00210755,0.00284838) (0.00967888,-0.0007969) (-0.00891201,-0.0163577) (-0.025356,-0.0138126) (0.00969038,0.0272957) (-0.0264836,0.0905323) (-0.00659636,-0.01184) (0.0779887,0.133857) (-0.132782,0.0892913) (0.0602514,-0.0141954) (-0.00468577,0.201334) (-0.00584357,0.0583142) (0.14252,0.182342) (-0.0680136,-0.0558422) (-0.0806263,-0.069619) (0.0693764,0.0172683) (-0.012331,0.0127468) (-0.00651142,-0.00190991) (0.00598103,-0.0043105) (-0.00079131,0.00044473) (-0.000517112,0.000835154) (0.000152274,-1.37794e-05) (3.42339e-05,-5.77791e-05) (-1.05241e-05,-3.17006e-06) (-1.68284e-06,2.09049e-06) (4.15773e-07,2.54252e-07) (5.76236e-08,-4.8373e-08) (-1.16341e-08,-9.56844e-09) (-1.21851e-09,8.98736e-10) (2.75589e-10,2.20068e-10) (1.27907e-11,-1.47704e-11) (-5.58138e-12,-3.2372e-12) (3.52389e-14,2.73991e-13) (1.13544e-13,2.0913e-14) (-8.72535e-15,-5.48044e-15) (-1.93234e-15,-2.18224e-16) (3.57439e-16,1.00058e-16) (2.37201e-17,1.48219e-17) (-8.4196e-18,-1.40488e-18) (-2.07791e-19,-4.30975e-19) 
  (5.93225e-24,-1.03266e-25) (-6.56228e-24,-6.98485e-23) (-9.00947e-22,6.88255e-23) (1.44734e-21,9.88812e-21) (1.18142e-19,-1.50005e-20) (-2.24094e-19,-1.21097e-18) (-1.3256e-17,2.21996e-18) (2.56843e-17,1.2735e-16) (1.26172e-15,-2.46435e-16) (-2.15277e-15,-1.13976e-14) (-1.00883e-13,2.09262e-14) (1.22039e-13,8.57861e-13) (6.69446e-12,-1.34525e-12) (-3.31236e-12,-5.33677e-11) (-3.62719e-10,6.28648e-11) (-1.27067e-10,2.67543e-09) (1.5679e-08,-1.89473e-09) (1.90019e-08,-1.04396e-07) (-5.23314e-07,1.95332e-08) (-1.03315e-06,3.03014e-06) (1.28709e-05,1.05323e-06) (3.24521e-05,-6.14232e-05) (-0.000216599,-4.91911e-05) (-0.000593107,0.000780031) (0.00218555,0.000811373) (0.0056018,-0.00496043) (-0.0104656,-0.00463135) (-0.0224012,0.00419618) (0.0121824,0.00389983) (0.03406,0.0604172) (-0.0184968,0.00701114) (0.10448,0.0152487) (-0.0124067,0.121981) (0.0100824,-0.0394693) (0.0991587,0.0968478) (0.0215225,0.0269619) (0.175399,0.0253563) (-0.0413004,0.00984444) (-0.0867507,0.0037338) (0.0397703,-0.024098) (0.00295122,0.0104858) (-0.00450193,0.00284781) (0.000679784,-0.00488353) (-0.00015848,0.000357165) (0.000160021,0.000692212) (8.28075e-05,-5.75371e-05) (-1.05751e-05,-4.96267e-05) (-7.94376e-06,2.14224e-06) (3.35261e-08,2.11525e-06) (3.72737e-07,-1.75937e-08) (1.39843e-08,-6.11003e-08) (-1.13511e-08,-8.27458e-10) (-4.64664e-10,1.26418e-09) (2.60148e-10,9.47331e-12) (5.69926e-12,-1.84678e-11) (-4.62807e-12,7.24356e-13) (5.17985e-14,2.15598e-13) (7.22523e-14,-4.41524e-14) (-6.07286e-15,-4.10833e-16) (-1.20085e-15,9.69773e-16) (2.16907e-16,-9.43107e-17) (2.20516e-17,-9.88956e-18) (-4.59676e-18,3.11652e-18) (-3.65887e-19,1.80899e-20) 
  (3.89476e-24,-2.45306e-24) (-3.07127e-23,-4.51557e-23) (-5.63062e-22,4.02213e-22) (4.65618e-21,6.08791e-21) (7.05519e-20,-5.57069e-20) (-5.96491e-19,-7.13194e-19) (-7.60972e-18,6.45291e-18) (6.37775e-17,7.25691e-17) (7.01777e-16,-6.18523e-16) (-5.61074e-15,-6.40164e-15) (-5.48933e-14,4.84403e-14) (3.99212e-13,4.86042e-13) (3.60069e-12,-3.05307e-12) (-2.24541e-11,-3.1218e-11) (-1.94779e-10,1.51864e-10) (9.65134e-10,1.64703e-09) (8.49498e-09,-5.79017e-09) (-3.00092e-08,-6.85982e-08) (-2.90097e-07,1.61499e-07) (6.11348e-07,2.14915e-06) (7.42158e-06,-3.07245e-06) (-6.40816e-06,-4.75147e-05) (-0.00013082,3.65101e-05) (-6.94687e-06,0.000668594) (0.00135758,-0.000248722) (0.000893796,-0.00497928) (-0.0059603,0.00116073) (-0.00955436,0.0122142) (0.00179174,-0.00312952) (0.0430868,0.0107114) (-0.00399,0.0202994) (0.0460716,-0.0438431) (0.0581426,0.0599776) (-0.0186887,-0.016894) (0.0850899,-0.00282626) (0.0158375,0.00206968) (0.0960833,-0.0704834) (-0.00151896,0.0149501) (-0.0422039,0.043822) (0.00565007,-0.0255313) (0.00637163,0.00140435) (-0.000617429,0.00350979) (-0.00183452,-0.00227541) (-1.47199e-05,0.000117289) (0.000382601,0.000239596) (2.88785e-05,-5.74242e-05) (-2.72678e-05,-1.95863e-05) (-3.83023e-06,4.26252e-06) (9.42268e-07,1.11856e-06) (2.07443e-07,-1.57911e-07) (-1.8796e-08,-4.17074e-08) (-6.72159e-09,3.95993e-09) (2.66985e-10,1.00463e-09) (1.45106e-10,-9.35159e-11) (-3.93269e-12,-1.59068e-11) (-2.0975e-12,2.13453e-12) (1.05526e-13,1.63276e-13) (1.69908e-14,-5.09171e-14) (-3.26297e-15,1.10148e-15) (-1.37977e-16,1.04985e-15) (6.58819e-17,-1.16368e-16) (4.75571e-18,-1.7644e-17) (-7.64337e-19,3.0792e-18) (-1.2381e-19,2.44788e-19) 
  (1.47176e-24,-2.87867e-24) (-3.48804e-23,-1.71426e-23) (-1.92839e-22,4.3961e-22) (4.94583e-21,2.08395e-21) (2.19866e-20,-5.74898e-20) (-6.00153e-19,-2.20003e-19) (-2.20178e-18,6.36773e-18) (6.18169e-17,2.05305e-17) (1.95779e-16,-5.90657e-16) (-5.35568e-15,-1.7327e-15) (-1.55259e-14,4.5313e-14) (3.86011e-13,1.33497e-13) (1.08244e-12,-2.83351e-12) (-2.27915e-11,-9.17801e-12) (-6.40739e-11,1.41832e-10) (1.07699e-09,5.3514e-10) (3.08426e-09,-5.55086e-09) (-3.93866e-08,-2.49258e-08) (-1.15632e-07,1.64834e-07) (1.06698e-06,8.72279e-07) (3.19264e-06,-3.57617e-06) (-2.02193e-05,-2.12952e-05) (-5.86632e-05,5.34149e-05) (0.000242697,0.000326341) (0.000599998,-0.000483565) (-0.00148773,-0.00266558) (-0.00217075,0.00190761) (0.000797064,0.00925194) (-0.00258377,0.000519549) (0.0209869,-0.0139931) (0.011222,0.0127297) (-0.00368688,-0.0343517) (0.0515018,-0.00324685) (-0.0140313,0.00468689) (0.032452,-0.0350348) (0.00431602,-0.00281909) (0.0106925,-0.071059) (0.00778153,-0.00229781) (-2.2516e-05,0.0376413) (-0.0074938,-0.0105158) (0.00261868,-0.00287986) (0.00127231,0.00166147) (-0.0015675,-0.000104374) (-3.94337e-05,5.22182e-05) (0.00025104,-5.79163e-05) (-2.45757e-06,-4.02159e-05) (-1.98259e-05,2.12326e-06) (-4.65361e-07,3.69567e-06) (8.94555e-07,1.78797e-07) (5.02363e-08,-1.60529e-07) (-2.64029e-08,-1.44602e-08) (-2.09267e-09,4.48285e-09) (5.53878e-10,4.53357e-10) (4.24453e-11,-9.68494e-11) (-8.95223e-12,-8.06431e-12) (-3.15178e-13,1.70652e-12) (1.3363e-13,7.11705e-14) (-1.01501e-14,-2.83545e-14) (-1.55886e-15,1.27813e-15) (3.67212e-16,5.30022e-16) (-6.05888e-18,-6.88152e-17) (-6.54784e-18,-1.03165e-17) (7.08142e-19,1.45939e-18) (8.67658e-20,1.67959e-19) 
  (-1.21831e-25,-2.09332e-24) (-2.54353e-23,1.77915e-24) (3.6708e-23,3.05139e-22) (3.43597e-21,-4.4549e-22) (-6.5713e-21,-3.83251e-20) (-3.98534e-19,7.1604e-20) (8.44269e-19,4.11554e-18) (3.94873e-17,-8.47182e-18) (-8.06951e-17,-3.74556e-16) (-3.32498e-15,7.58545e-16) (5.6479e-15,2.85937e-14) (2.36321e-13,-5.09487e-14) (-2.69921e-13,-1.80595e-12) (-1.40126e-11,2.45617e-12) (6.75947e-12,9.25713e-11) (6.79181e-10,-7.39136e-11) (1.05639e-10,-3.7559e-09) (-2.6093e-08,5.11498e-10) (-1.74403e-08,1.17086e-07) (7.62049e-07,6.53458e-08) (7.43427e-07,-2.69619e-06) (-1.59297e-05,-3.06331e-06) (-1.61175e-05,4.24573e-05) (0.000215005,6.15833e-05) (0.00016852,-0.000386353) (-0.00155589,-0.000591217) (-0.000556478,0.00120873) (0.00375928,0.00324377) (-0.000558989,0.00289158) (0.0016499,-0.0127735) (0.0117921,-0.000392807) (-0.0148402,-0.0086877) (0.0177747,-0.0232805) (-0.00188836,0.00798065) (-0.000621263,-0.0248924) (0.000636064,-0.000200385) (-0.0239032,-0.0313659) (-0.000547125,-0.00837566) (0.0145623,0.0150298) (-0.00563967,-0.000384201) (-0.000541467,-0.00217428) (0.00109714,9.58164e-05) (-0.000559939,0.000540585) (-2.26116e-05,6.30422e-05) (7.0791e-05,-0.000113864) (-1.4642e-05,-1.94745e-05) (-7.33235e-06,7.95899e-06) (1.1066e-06,1.96419e-06) (4.68396e-07,-2.35422e-07) (-3.24526e-08,-9.54874e-08) (-1.8035e-08,2.59781e-09) (4.85365e-10,2.89581e-09) (4.48229e-10,2.471e-11) (-9.46173e-12,-6.02923e-11) (-7.83443e-12,-9.20064e-13) (3.36278e-13,8.7856e-13) (1.02326e-13,-9.00872e-15) (-1.2535e-14,-8.6398e-15) (-5.39074e-16,1.07234e-15) (3.44222e-16,8.73827e-17) (-2.02375e-17,-2.67702e-17) (-7.18357e-18,-1.55137e-18) (6.71663e-19,3.43516e-19) (1.15086e-19,2.59211e-20) 
  (-7.04373e-25,-1.05857e-24) (-1.28072e-23,8.81776e-24) (1.11472e-22,1.46114e-22) (1.64029e-21,-1.28006e-21) (-1.48505e-20,-1.74521e-20) (-1.80878e-19,1.5588e-19) (1.64613e-18,1.80297e-18) (1.71432e-17,-1.57987e-17) (-1.49892e-16,-1.60827e-16) (-1.3952e-15,1.32121e-15) (1.1041e-14,1.23288e-14) (9.71992e-14,-9.0328e-14) (-6.45058e-13,-8.02163e-13) (-5.74067e-12,4.98947e-12) (2.90849e-11,4.32766e-11) (2.81917e-10,-2.18525e-10) (-9.72618e-10,-1.87448e-09) (-1.11707e-08,7.36918e-09) (2.2836e-08,6.2732e-08) (3.41501e-07,-1.84684e-07) (-3.55064e-07,-1.5388e-06) (-7.48985e-06,3.33031e-06) (3.53121e-06,2.51268e-05) (0.000104921,-4.05414e-05) (-2.06139e-05,-0.000227445) (-0.000779664,0.000277452) (-4.97001e-05,0.000658793) (0.0023851,-0.000198469) (0.00150522,0.00169924) (-0.00409633,-0.00433596) (0.00450734,-0.00566716) (-0.00724397,0.00330659) (-0.00298697,-0.0151277) (0.00287617,0.00314174) (-0.00860208,-0.00872459) (0.00122272,0.000546245) (-0.019795,-0.0021194) (-0.00577281,-0.00348868) (0.0105752,0.000286525) (-0.00138681,0.00173863) (-0.00110447,-0.00047928) (0.00038566,-0.000360354) (1.39601e-05,0.000359689) (1.55207e-05,4.80643e-05) (-1.4826e-05,-6.25813e-05) (-1.33435e-05,-3.93818e-06) (-1.971e-07,5.4408e-06) (1.17338e-06,4.87172e-07) (1.22816e-07,-2.53912e-07) (-4.6593e-08,-3.19167e-08) (-7.26883e-09,7.28211e-09) (1.14682e-09,1.17674e-09) (2.18082e-10,-1.42297e-10) (-2.20813e-11,-2.53676e-11) (-4.10911e-12,2.27792e-12) (3.76453e-13,3.14754e-13) (4.79155e-14,-3.9429e-14) (-7.0545e-15,-2.4578e-16) (1.93135e-17,6.82299e-16) (1.61492e-16,-7.80378e-17) (-1.45268e-17,-6.12052e-18) (-3.4304e-18,2.12791e-18) (3.24368e-19,-3.47937e-20) (5.51847e-20,-3.8014e-20) 
  (-6.53202e-25,-3.18481e-25) (-3.70756e-24,8.07322e-24) (9.58598e-23,3.89638e-23) (4.23494e-22,-1.09214e-21) (-1.20137e-20,-4.10464e-21) (-4.18266e-20,1.25373e-19) (1.27524e-18,3.81622e-19) (3.62906e-18,-1.21174e-17) (-1.13596e-16,-3.23959e-17) (-2.82336e-16,9.78804e-16) (8.40356e-15,2.56945e-15) (1.98419e-14,-6.55995e-14) (-5.09323e-13,-1.86642e-13) (-1.23409e-12,3.61589e-12) (2.48021e-11,1.16957e-11) (6.5228e-11,-1.61788e-10) (-9.45457e-10,-5.9105e-10) (-2.79525e-09,5.76346e-09) (2.74111e-08,2.26448e-08) (9.12989e-08,-1.59097e-07) (-5.85697e-07,-6.1236e-07) (-2.05981e-06,3.2449e-06) (8.6055e-06,1.05174e-05) (2.80625e-05,-4.41117e-05) (-7.18145e-05,-9.70339e-05) (-0.000188652,0.000327286) (0.000122555,0.000336004) (0.0006484,-0.000820538) (0.00141894,-2.35703e-05) (-0.00251226,0.000297237) (-0.000741575,-0.00394907) (-0.000542007,0.00345041) (-0.00651169,-0.00388567) (0.00205364,-0.000217157) (-0.00575602,-0.000320244) (0.00124757,-0.000384517) (-0.00701011,0.00614381) (-0.00420373,0.00140513) (0.00358246,-0.00334302) (0.000345162,0.000752261) (-0.000533196,0.000264129) (-7.72452e-06,-0.00023349) (0.000121586,9.9236e-05) (2.72098e-05,1.54321e-05) (-2.44438e-05,-1.49529e-05) (-6.85756e-06,2.86074e-06) (1.57487e-06,2.03148e-06) (6.40611e-07,-1.9101e-07) (-2.84408e-08,-1.4098e-07) (-2.96568e-08,1.49354e-09) (-7.64894e-10,5.42015e-09) (8.56633e-10,1.62279e-10) (4.95927e-11,-1.3232e-10) (-1.70616e-11,-5.1629e-12) (-1.1066e-12,2.33953e-12) (2.46457e-13,5.2332e-14) (9.39641e-15,-3.27842e-14) (-2.75584e-15,1.37623e-15) (1.93774e-16,3.00846e-16) (3.5514e-17,-7.6017e-17) (-7.25395e-18,8.15786e-19) (-5.3764e-19,1.97831e-18) (1.12433e-19,-7.75208e-20) (6.13745e-21,-3.44625e-20) 
  (-3.92409e-25,3.11187e-26) (5.24447e-25,4.75905e-24) (5.4567e-23,-8.21077e-24) (-1.06524e-22,-6.13021e-22) (-6.50777e-21,1.38189e-21) (1.50544e-20,6.74249e-20) (6.63489e-19,-1.70203e-19) (-1.5926e-18,-6.29442e-18) (-5.7605e-17,1.57853e-17) (1.27782e-16,4.95964e-16) (4.23955e-15,-1.08847e-15) (-7.69849e-15,-3.27663e-14) (-2.62147e-13,5.27225e-14) (3.38012e-13,1.79753e-12) (1.33861e-11,-1.47382e-12) (-1.00465e-11,-8.07576e-11) (-5.49858e-10,-4.20931e-12) (1.60961e-10,2.91808e-09) (1.75632e-08,2.38066e-09) (-6.37566e-11,-8.23516e-08) (-4.14827e-07,-1.01327e-07) (-1.28932e-08,1.70087e-06) (6.56787e-06,2.0359e-06) (-1.10601e-06,-2.26871e-05) (-5.75296e-05,-2.02728e-05) (2.81486e-05,0.000156602) (0.000150673,0.000120263) (-7.46291e-05,-0.00040843) (0.000499073,-0.000586646) (-0.000436915,0.000900184) (-0.00176524,-0.00103855) (0.00112375,0.000968191) (-0.00335646,0.00100244) (0.000501411,-0.000789039) (-0.00205465,0.00162859) (0.000394307,-0.000804846) (-4.07342e-05,0.00407476) (-0.00102246,0.00232293) (7.95331e-05,-0.00208695) (0.000333257,-3.55003e-05) (-7.32201e-05,0.000259446) (-7.61171e-05,-5.99316e-05) (6.40863e-05,-1.07588e-05) (1.64642e-05,-4.36346e-06) (-1.15811e-05,2.82947e-06) (-1.65475e-06,3.31988e-06) (1.12178e-06,2.60844e-07) (1.82004e-07,-2.7507e-07) (-5.25685e-08,-4.63576e-08) (-1.12141e-08,9.56849e-09) (1.34091e-09,2.41494e-09) (4.0084e-10,-1.83202e-10) (-1.97047e-11,-6.96258e-11) (-8.77485e-12,2.46035e-12) (2.35467e-13,1.31464e-12) (1.23381e-13,-3.54448e-14) (-5.38483e-15,-1.65064e-14) (-8.38341e-16,1.01935e-15) (1.55423e-16,7.21159e-17) (-8.49242e-18,-3.5616e-17) (-2.69295e-18,1.97901e-18) (4.41762e-19,8.65893e-19) (3.02247e-20,-5.04791e-20) (-9.4448e-21,-1.41174e-20) 
  (-1.65674e-25,1.17187e-25) (1.48628e-24,1.94519e-24) (2.16278e-23,-1.77811e-23) (-2.06054e-22,-2.36185e-22) (-2.42473e-21,2.25969e-21) (2.3741e-20,2.46933e-20) (2.34388e-19,-2.38653e-19) (-2.25192e-18,-2.22402e-18) (-1.96372e-17,2.07623e-17) (1.74067e-16,1.7261e-16) (1.43242e-15,-1.47348e-15) (-1.08509e-14,-1.14858e-14) (-9.06122e-14,8.42402e-14) (5.39955e-13,6.4556e-13) (4.87746e-12,-3.806e-12) (-2.12721e-11,-2.99372e-11) (-2.15971e-10,1.32325e-10) (6.6564e-10,1.11257e-09) (7.49392e-09,-3.46541e-09) (-1.70255e-08,-3.16552e-08) (-1.89354e-07,6.86771e-08) (3.60062e-07,6.297e-07) (3.11e-06,-1.00073e-06) (-5.56099e-06,-7.52537e-06) (-2.7838e-05,8.47327e-06) (4.72503e-05,4.0271e-05) (9.74816e-05,3.10544e-06) (-0.000131646,-7.13262e-05) (-5.42306e-05,-0.000370856) (0.00023132,0.000308636) (-0.000920632,0.000304771) (0.000591505,-0.000196899) (-0.000681358,0.0013668) (-0.000116537,-0.000378878) (-0.000205357,0.00114208) (-0.000197862,-0.000477192) (0.00125484,0.00110622) (0.000516733,0.00120331) (-0.000557762,-0.000600955) (3.95268e-05,-0.000156446) (5.72218e-05,9.62458e-05) (-3.73069e-05,8.51373e-06) (1.34809e-05,-2.1856e-05) (4.20023e-06,-7.3175e-06) (-2.40608e-06,3.97522e-06) (4.67883e-07,1.67244e-06) (4.4708e-07,-2.12074e-07) (-1.8429e-08,-1.52259e-07) (-3.27325e-08,-2.29038e-09) (-1.41916e-09,6.80317e-09) (1.2167e-09,5.33072e-10) (1.06115e-10,-1.84822e-10) (-2.77999e-11,-2.15973e-11) (-2.9641e-12,3.38006e-12) (4.63908e-13,4.58688e-13) (4.54618e-14,-4.5739e-14) (-6.4899e-15,-5.20174e-15) (-1.85866e-16,5.53686e-16) (7.44105e-17,-9.33739e-18) (-1.16856e-17,-9.34811e-18) (-5.64892e-19,1.38581e-18) (4.0419e-19,1.57511e-19) (3.11514e-21,-2.69041e-20) (-7.5095e-21,-1.80913e-21) 
  (-4.02362e-26,9.14405e-26) (1.11097e-24,4.35175e-25) (4.52344e-24,-1.27901e-23) (-1.4344e-22,-4.51626e-23) (-4.30237e-22,1.51658e-21) (1.56449e-20,4.07447e-21) (3.57166e-20,-1.51639e-19) (-1.43003e-18,-3.34652e-19) (-2.73912e-18,1.27189e-17) (1.08708e-16,2.63089e-17) (2.04816e-16,-8.91475e-16) (-6.81628e-15,-1.97246e-15) (-1.4739e-14,5.19791e-14) (3.49036e-13,1.31445e-13) (9.44309e-13,-2.49916e-12) (-1.44468e-11,-7.16703e-12) (-4.94028e-11,9.76462e-11) (4.81046e-10,2.98419e-10) (1.94433e-09,-3.03733e-09) (-1.28276e-08,-8.75726e-09) (-5.23048e-08,7.21338e-08) (2.60056e-07,1.58582e-07) (8.59471e-07,-1.17661e-06) (-3.46221e-06,-1.37475e-06) (-7.50278e-06,1.06769e-05) (2.2523e-05,1.00492e-06) (3.57663e-05,-2.83653e-05) (-4.38117e-05,2.21947e-05) (-0.000140503,-8.93863e-05) (0.000151632,-3.81483e-05) (-0.000167575,0.000396205) (5.79043e-05,-0.000255904) (0.000213336,0.000593803) (-0.000142856,-6.82262e-05) (0.000261851,0.000427065) (-0.000253012,-8.0927e-05) (0.000640528,-0.000100623) (0.000583085,0.000213205) (-0.000295366,-9.19202e-06) (-5.92071e-05,-5.60242e-05) (4.13606e-05,1.02293e-05) (-6.21605e-06,1.3284e-05) (-2.85182e-06,-9.28244e-06) (-1.06408e-06,-3.72864e-06) (4.02489e-07,1.65021e-06) (6.54086e-07,3.98309e-07) (9.21857e-08,-1.8391e-07) (-4.98605e-08,-4.5569e-08) (-1.22914e-08,8.23291e-09) (1.37291e-09,2.81142e-09) (5.92995e-10,-1.46636e-10) (-1.03644e-11,-9.83968e-11) (-1.63549e-11,-4.2304e-13) (-2.78852e-13,2.12063e-12) (2.99764e-13,5.18497e-14) (7.73914e-15,-3.06123e-14) (-3.77925e-15,-4.28317e-16) (1.1676e-17,2.71844e-16) (2.39451e-17,-1.83489e-17) (-5.72818e-18,-9.98941e-20) (1.2659e-19,6.34027e-19) (1.72337e-19,-6.27262e-20) (-4.68403e-21,-1.20634e-20) (-2.92847e-21,1.56062e-21) 
  (6.12481e-27,4.67018e-26) (5.48198e-25,-9.64576e-26) (-1.2961e-24,-6.16081e-24) (-6.68964e-23,1.6818e-23) (1.92892e-22,6.91746e-22) (6.96079e-21,-2.14781e-21) (-2.16266e-20,-6.60143e-20) (-6.16003e-19,2.07161e-19) (1.85425e-18,5.35162e-18) (4.62926e-17,-1.49632e-17) (-1.20588e-16,-3.69102e-16) (-2.94302e-15,7.75677e-16) (5.77076e-15,2.16645e-14) (1.56682e-13,-2.55008e-14) (-1.87249e-13,-1.07634e-12) (-6.8695e-12,2.71075e-13) (3.12077e-12,4.45801e-11) (2.42679e-10,1.71859e-11) (1.65883e-11,-1.48727e-09) (-6.63359e-09,-7.6173e-10) (-1.25441e-09,3.71314e-08) (1.27514e-07,6.183e-09) (-3.20184e-09,-6.11703e-07) (-1.44758e-06,2.22961e-07) (3.80869e-07,5.48865e-06) (6.46645e-06,-4.16709e-06) (3.12787e-06,-1.95605e-05) (-1.77932e-07,1.49783e-05) (-6.51404e-05,2.07463e-05) (1.09839e-05,-6.86378e-05) (7.84724e-05,0.000161969) (-7.70885e-05,-7.85803e-05) (0.000225389,0.000103392) (-5.67409e-05,1.99155e-05) (0.000202369,5.83708e-05) (-0.000105496,6.81592e-05) (0.000117096,-0.000208014) (0.000245077,-0.000122076) (-6.96298e-05,6.72342e-05) (-3.82186e-05,6.99553e-06) (1.27529e-05,-7.48937e-06) (2.54772e-06,4.92965e-06) (-3.20542e-06,-1.44586e-06) (-1.47746e-06,-7.86398e-07) (4.94567e-07,3.05887e-07) (3.12035e-07,-6.83943e-08) (-1.61969e-08,-8.1735e-08) (-2.83021e-08,-8.03705e-10) (-1.97003e-09,6.12031e-09) (1.21399e-09,5.95483e-10) (1.67024e-10,-2.11335e-10) (-2.97142e-11,-3.27605e-11) (-5.98475e-12,4.17379e-12) (4.44211e-13,8.74828e-13) (1.23801e-13,-5.71875e-14) (-4.57124e-15,-1.42199e-14) (-1.526e-15,7.08229e-16) (5.71187e-17,1.16486e-16) (4.92207e-18,-1.01842e-17) (-1.63752e-18,1.22238e-18) (1.9417e-19,1.82971e-19) (3.57486e-20,-6.46468e-20) (-4.89083e-21,-3.64716e-21) (-4.93752e-22,1.26354e-21) 
  (1.34023e-26,1.65857e-26) (1.86735e-25,-1.65305e-25) (-1.93138e-24,-2.03401e-24) (-2.11312e-23,2.17855e-23) (2.30786e-22,2.13038e-22) (2.05838e-21,-2.37524e-21) (-2.2706e-20,-1.92023e-20) (-1.74482e-19,2.12278e-19) (1.82513e-18,1.50542e-18) (1.30473e-17,-1.53937e-17) (-1.19155e-16,-1.03744e-16) (-8.64221e-16,8.95003e-16) (6.30219e-15,6.28772e-15) (4.98417e-14,-4.11081e-14) (-2.70973e-13,-3.30087e-13) (-2.41094e-12,1.47612e-12) (9.64816e-12,1.45311e-11) (9.27299e-11,-4.25821e-11) (-2.95254e-10,-5.05289e-10) (-2.61689e-09,1.08143e-09) (7.68656e-09,1.25447e-08) (4.76357e-08,-2.40026e-08) (-1.45218e-07,-1.94608e-07) (-4.50883e-07,3.61546e-07) (1.50941e-06,1.58032e-06) (1.09635e-06,-2.27724e-06) (-4.59536e-06,-6.56813e-06) (4.46765e-06,1.45091e-06) (-9.30785e-06,2.44742e-05) (-2.57081e-05,-1.9463e-05) (6.88632e-05,1.88781e-05) (-4.4783e-05,7.33564e-06) (8.73167e-05,-3.21882e-05) (-1.06101e-05,1.93826e-05) (7.64311e-05,-3.93144e-05) (-5.64358e-06,5.53317e-05) (-3.41197e-05,-7.68717e-05) (3.30355e-05,-0.000108358) (2.52662e-07,2.8124e-05) (-8.49238e-06,1.47841e-05) (1.3179e-06,-4.43923e-06) (2.05438e-06,3.97994e-07) (-1.11005e-06,5.01861e-07) (-6.50086e-07,2.13206e-07) (1.8132e-07,-3.93427e-08) (6.96837e-08,-1.05596e-07) (-2.49937e-08,-2.15549e-08) (-8.79612e-09,7.16904e-09) (9.68206e-10,2.51445e-09) (5.51733e-10,-1.14881e-10) (6.39722e-13,-1.14192e-10) (-1.87141e-11,-3.72431e-12) (-1.00555e-12,2.96936e-12) (3.82945e-13,2.04323e-13) (3.02225e-14,-5.07806e-14) (-5.27622e-15,-4.28857e-15) (-4.10096e-16,6.00795e-16) (4.85722e-17,3.69819e-17) (3.4073e-19,-4.10637e-18) (-1.71821e-19,6.46718e-19) (1.04006e-19,1.09119e-20) (-5.94576e-21,-2.78681e-20) (-2.75817e-21,-6.49371e-23) (1.67028e-22,5.04607e-22) 
  (8.76716e-27,3.0781e-27) (3.1005e-26,-1.03065e-25) (-1.16365e-24,-3.02162e-25) (-2.70795e-24,1.25601e-23) (1.29826e-22,2.44664e-23) (1.98775e-22,-1.28702e-21) (-1.21133e-20,-1.7569e-21) (-1.40113e-20,1.10363e-19) (9.41032e-19,1.30763e-19) (1.15333e-18,-7.90313e-18) (-6.08146e-17,-1.09677e-17) (-1.05758e-16,4.72362e-16) (3.28105e-15,8.99458e-16) (8.60387e-15,-2.3532e-14) (-1.49244e-13,-6.105e-14) (-5.39662e-13,9.75583e-13) (5.81161e-12,3.12833e-12) (2.41517e-11,-3.35977e-11) (-1.92735e-10,-1.11607e-10) (-7.05263e-10,9.32595e-10) (5.02273e-09,2.45e-09) (1.16786e-08,-1.85874e-08) (-8.75441e-08,-2.71736e-08) (-8.00095e-08,2.14703e-07) (8.14952e-07,9.03202e-08) (-1.97915e-08,-8.42244e-07) (-2.99802e-06,-5.1781e-07) (9.07258e-07,-1.52473e-06) (5.10414e-06,7.96452e-06) (-1.37605e-05,4.97754e-06) (2.24945e-05,-1.49103e-05) (-8.58736e-06,1.59659e-05) (1.45029e-05,-3.01853e-05) (1.44615e-06,7.93554e-06) (1.07528e-05,-3.21766e-05) (1.68185e-05,1.62127e-05) (-2.81266e-05,-5.43363e-06) (-2.19092e-05,-3.84355e-05) (5.12798e-06,4.49098e-06) (2.0706e-06,6.58317e-06) (-5.27186e-07,-1.16067e-06) (6.10483e-07,-4.94988e-07) (-1.17002e-07,3.85513e-07) (-1.15084e-07,2.40179e-07) (3.11757e-08,-4.48081e-08) (-9.27195e-09,-4.68153e-08) (-1.27836e-08,-5.01505e-10) (-7.64771e-10,4.30013e-09) (9.47827e-10,5.3636e-10) (1.46908e-10,-1.73549e-10) (-2.86256e-11,-3.68424e-11) (-7.17539e-12,3.44296e-12) (3.96747e-13,1.24017e-12) (1.83783e-13,-2.39141e-14) (-1.58259e-15,-2.48058e-14) (-2.96474e-15,-2.73487e-16) (-1.97082e-17,3.08782e-16) (2.75148e-17,4.12436e-18) (-2.91854e-19,-1.56555e-18) (8.32554e-20,1.75761e-19) (3.24472e-20,-2.1367e-20) (-8.46247e-21,-6.34664e-21) (-9.56899e-22,7.02538e-22) (1.68789e-22,1.09217e-22) 
  (3.81175e-27,-8.52958e-28) (-1.17919e-26,-4.32673e-26) (-4.73312e-25,1.50731e-25) (1.79784e-24,4.92956e-24) (4.97223e-23,-1.98044e-23) (-2.07812e-22,-4.76179e-22) (-4.42534e-21,1.98014e-21) (1.8356e-20,3.91381e-20) (3.35039e-19,-1.49455e-19) (-1.21677e-18,-2.76424e-18) (-2.17451e-17,8.21908e-18) (5.73025e-17,1.69763e-16) (1.21866e-15,-3.00704e-16) (-1.61135e-15,-9.10451e-15) (-5.9123e-14,5.28858e-15) (3.86647e-15,4.20761e-13) (2.45688e-12,6.11217e-14) (1.56242e-12,-1.60608e-11) (-8.32174e-11,-2.39691e-12) (-4.4441e-11,4.63606e-10) (2.05209e-09,-1.94553e-10) (-9.37125e-11,-8.7813e-09) (-3.15216e-08,1.02692e-08) (1.89703e-08,8.81413e-08) (2.42783e-07,-1.61225e-07) (-1.34575e-07,-2.71223e-07) (-8.76825e-07,6.44393e-07) (-4.87089e-07,-5.88912e-07) (3.27725e-06,7.24442e-08) (-1.79756e-06,6.04945e-06) (1.28368e-06,-9.6703e-06) (2.60123e-06,6.45489e-06) (-3.51388e-06,-1.10664e-05) (2.21815e-06,2.03924e-06) (-5.82496e-06,-1.1532e-05) (9.29154e-06,-1.35997e-06) (-6.63303e-06,6.88178e-06) (-1.59265e-05,-3.83999e-06) (1.07469e-06,-2.85226e-07) (2.31204e-06,1.17176e-06) (-2.52693e-07,-1.43288e-07) (1.65092e-08,-2.91506e-07) (6.81913e-08,1.06909e-07) (3.49687e-08,9.27422e-08) (-1.50424e-09,-1.44228e-08) (-1.4279e-08,-9.57043e-09) (-3.86863e-09,2.91805e-09) (8.23531e-10,1.39649e-09) (4.1782e-10,-7.67106e-11) (3.23851e-12,-8.90022e-11) (-1.78813e-11,-4.41128e-12) (-1.46542e-12,2.86023e-12) (4.25597e-13,3.06156e-13) (5.56411e-14,-5.2471e-14) (-6.28682e-15,-8.003e-15) (-1.09786e-15,6.106e-16) (5.95642e-17,1.15172e-16) (1.13656e-17,-4.5071e-18) (-3.0135e-19,-6.28725e-19) (4.38113e-20,1.46647e-20) (3.48832e-21,-1.32411e-20) (-3.78666e-21,2.98811e-22) (-1.21926e-22,4.70977e-22) (7.36424e-23,-6.57621e-24) 
  (1.12593e-27,-1.11915e-27) (-1.33328e-26,-1.22064e-26) (-1.26915e-25,1.52267e-25) (1.64443e-24,1.25968e-24) (1.21505e-23,-1.70202e-23) (-1.66273e-22,-1.11204e-22) (-1.0096e-21,1.54869e-21) (1.36575e-20,8.63063e-21) (7.52706e-20,-1.13382e-19) (-9.04119e-19,-6.13355e-19) (-5.18568e-18,6.60065e-18) (4.80315e-17,4.09465e-17) (3.28247e-16,-3.03431e-16) (-2.06157e-15,-2.51321e-15) (-1.82228e-14,1.12768e-14) (7.46751e-14,1.3278e-13) (8.26317e-13,-3.81567e-13) (-2.52253e-12,-5.50097e-12) (-2.77878e-11,1.3628e-11) (8.05251e-11,1.5902e-10) (6.05701e-10,-4.38702e-10) (-1.92596e-09,-2.78499e-09) (-7.08e-09,9.18244e-09) (2.52184e-08,2.38042e-08) (2.87111e-08,-9.41679e-08) (-9.50516e-08,-6.88195e-08) (-4.42495e-08,3.65363e-07) (-3.15254e-07,7.05359e-08) (5.97437e-07,-9.46727e-07) (1.46804e-06,2.11008e-06) (-2.23464e-06,-2.54089e-06) (2.4081e-06,8.65012e-07) (-3.3798e-06,-1.94633e-06) (1.16146e-06,1.10349e-07) (-4.53317e-06,-1.38604e-06) (1.7723e-06,-3.17451e-06) (7.97981e-07,3.06724e-06) (-4.82062e-06,3.17411e-06) (-1.75376e-07,-1.77049e-08) (8.66419e-07,-2.713e-07) (-4.752e-08,-1.16115e-08) (-7.14871e-08,-7.90333e-08) (3.76345e-08,4.37076e-09) (3.25303e-08,1.38512e-08) (-2.21115e-09,-2.50993e-09) (-5.80531e-09,1.17467e-09) (-3.97482e-10,1.74439e-09) (5.50966e-10,1.89659e-10) (1.01359e-10,-1.23872e-10) (-2.01028e-11,-2.73354e-11) (-6.40609e-12,2.92431e-12) (2.28057e-13,1.23706e-12) (2.05102e-13,-3.30305e-15) (5.53641e-15,-3.00445e-14) (-3.88233e-15,-1.19744e-15) (-2.26219e-16,4.59402e-16) (4.57918e-17,2.75131e-17) (3.14671e-18,-4.12901e-18) (-2.35846e-19,-2.27282e-19) (4.15159e-21,-6.91623e-21) (-2.34624e-21,-3.97252e-21) (-9.15398e-22,9.60932e-22) (8.30678e-23,1.71658e-22) (1.96214e-23,-1.79913e-23) 
  (1.37279e-28,-6.09877e-28) (-6.95618e-27,-1.20883e-27) (-9.28333e-27,7.5986e-26) (7.89327e-25,6.30618e-26) (3.26251e-25,-7.88592e-24) (-7.44441e-23,-9.59124e-25) (1.96848e-24,6.78949e-22) (5.81563e-21,-6.23985e-23) (6.02454e-22,-4.84187e-20) (-3.78082e-19,-1.33533e-20) (-3.41992e-19,2.87726e-18) (2.08341e-17,3.74443e-18) (4.91053e-17,-1.45073e-16) (-1.00906e-15,-4.21958e-16) (-4.03391e-15,6.43889e-15) (4.47129e-14,2.90388e-14) (2.1107e-13,-2.61343e-13) (-1.78335e-12,-1.27617e-12) (-6.74475e-12,9.3031e-12) (5.64817e-11,3.33577e-11) (1.09613e-10,-2.46239e-10) (-1.17511e-09,-4.37624e-10) (-2.98981e-10,3.95398e-09) (1.27934e-08,1.61772e-09) (-1.16903e-08,-2.95061e-08) (-4.6258e-08,-2.69146e-09) (7.62948e-08,8.99365e-08) (-3.89734e-08,1.216e-07) (-1.88692e-07,-3.40934e-07) (9.86597e-07,8.96351e-08) (-1.12953e-06,2.92194e-09) (8.04459e-07,-4.06492e-07) (-1.25047e-06,2.60087e-07) (3.84338e-07,-2.55933e-07) (-1.44974e-06,8.39166e-07) (-5.39905e-07,-1.24967e-06) (1.01433e-06,2.92486e-07) (-3.20986e-07,1.91259e-06) (-5.55229e-08,2.00905e-07) (1.47906e-07,-2.58236e-07) (-1.04351e-08,-1.19583e-08) (-3.79633e-08,-3.04446e-09) (7.33697e-09,-7.88471e-09) (1.1125e-08,-4.78148e-09) (-5.68888e-10,-3.34671e-10) (-1.06459e-09,1.63961e-09) (3.03433e-10,5.6619e-10) (1.89551e-10,-7.41555e-11) (-1.35425e-12,-5.83076e-11) (-1.21642e-11,-3.24477e-12) (-1.18632e-12,2.32974e-12) (3.5687e-13,3.17673e-13) (6.17898e-14,-4.78262e-14) (-5.19998e-15,-1.06305e-14) (-1.5065e-15,4.85308e-16) (3.07008e-17,1.99898e-16) (2.15573e-17,-5.4634e-19) (2.08608e-19,-2.12719e-18) (-1.44997e-19,-4.68661e-20) (-4.60734e-21,-5.56407e-22) (-1.50304e-21,-2.48309e-22) (-8.27038e-24,4.543e-22) (6.61726e-23,2.80355e-23) (1.70483e-24,-9.28515e-24) 
  (-8.21558e-29,-2.24415e-28) (-2.46103e-27,1.05141e-27) (1.26738e-26,2.57133e-26) (2.57285e-25,-1.41241e-25) (-1.49398e-24,-2.46481e-24) (-2.25416e-23,1.45306e-23) (1.34248e-22,1.99298e-22) (1.67286e-21,-1.12842e-21) (-8.90871e-21,-1.38774e-20) (-1.08234e-19,6.3093e-20) (3.9807e-19,8.63034e-19) (6.38369e-18,-2.21387e-18) (-8.03785e-18,-4.96011e-17) (-3.54936e-16,2.02563e-17) (-2.8907e-16,2.62712e-15) (1.81473e-14,2.18665e-15) (2.56947e-14,-1.2022e-13) (-7.69354e-13,-8.77362e-14) (-5.30702e-13,4.20706e-12) (2.32951e-11,-7.62995e-13) (-1.07213e-11,-9.61726e-11) (-4.31048e-10,1.14753e-10) (6.33643e-10,1.18134e-09) (3.98689e-09,-2.31307e-09) (-8.40672e-09,-5.09365e-09) (-1.48665e-08,9.80408e-09) (3.57692e-08,1.47836e-09) (3.1236e-08,3.57492e-08) (-1.40947e-07,7.34345e-10) (2.61433e-07,-2.51273e-07) (-2.39613e-07,2.73655e-07) (9.54394e-08,-2.89702e-07) (-2.47781e-07,3.27155e-07) (4.6204e-08,-1.76169e-07) (-1.19027e-07,5.57765e-07) (-4.78931e-07,-1.21277e-07) (2.58291e-07,-2.4187e-07) (3.81645e-07,4.91832e-07) (6.93842e-08,9.75674e-08) (-1.77787e-08,-8.97948e-08) (-8.44358e-09,-5.89879e-09) (-1.06289e-08,8.0256e-09) (-8.10291e-10,-2.86632e-09) (1.38338e-09,-3.73738e-09) (-1.4711e-10,-1.35997e-10) (1.37886e-10,6.0295e-10) (2.10483e-10,7.63422e-11) (3.29008e-11,-6.10245e-11) (-1.38271e-11,-1.52498e-11) (-4.15311e-12,1.8631e-12) (1.89606e-13,9.2539e-13) (1.75966e-13,1.08301e-14) (7.62539e-15,-2.79977e-14) (-3.96093e-15,-2.03617e-15) (-3.60595e-16,4.81929e-16) (5.37828e-17,5.59421e-17) (6.99086e-18,-4.83947e-18) (-3.84192e-19,-7.6501e-19) (-6.64692e-20,1.38723e-20) (-2.23467e-21,2.54334e-21) (-3.63235e-22,3.73693e-22) (1.03544e-22,1.13634e-22) (2.4758e-23,-8.51065e-24) (-1.48476e-24,-2.95958e-24) 
  (-7.11927e-29,-5.31725e-29) (-5.43652e-28,8.22498e-28) (9.01995e-27,5.23863e-27) (4.8579e-26,-9.37939e-26) (-9.27119e-25,-4.26021e-25) (-3.65732e-24,8.61455e-24) (7.6267e-23,3.01977e-23) (2.51652e-22,-6.25761e-22) (-4.92665e-21,-2.11479e-21) (-1.80634e-20,3.51574e-20) (2.44292e-19,1.62966e-19) (1.39461e-18,-1.49978e-18) (-9.19236e-18,-1.27553e-17) (-1.01272e-16,5.10771e-17) (2.92713e-16,8.53402e-16) (5.94148e-15,-1.91435e-15) (-1.18185e-14,-4.26916e-14) (-2.49857e-13,1.00297e-13) (5.93473e-13,1.42287e-12) (6.67589e-12,-4.49249e-12) (-2.10004e-11,-2.7329e-11) (-9.76069e-11,1.17568e-10) (3.92786e-10,2.2244e-10) (5.874e-10,-1.46745e-09) (-2.95087e-09,2.08486e-10) (-1.92218e-09,6.25442e-09) (7.30717e-09,-7.19623e-09) (1.66762e-08,-3.16174e-09) (-2.65042e-08,4.51443e-08) (-5.01716e-09,-1.26436e-07) (1.40714e-08,1.12337e-07) (-4.239e-08,-9.01723e-08) (8.43235e-09,1.29809e-07) (-3.42946e-08,-6.12812e-08) (1.11797e-07,1.50247e-07) (-1.37112e-07,1.07046e-07) (-2.35834e-08,-1.16186e-07) (1.90489e-07,1.52724e-08) (5.34973e-08,6.38585e-09) (-2.02309e-08,-1.71893e-08) (-4.95844e-09,-1.07402e-10) (-9.8211e-10,4.45137e-09) (-8.52413e-10,-1.32881e-10) (-5.59189e-10,-1.12987e-09) (-9.3678e-11,-5.26123e-11) (1.61013e-10,9.63079e-11) (6.98031e-11,-2.92458e-11) (-4.80153e-12,-2.25851e-11) (-7.00025e-12,-8.28332e-13) (-7.12246e-13,1.43754e-12) (2.55905e-13,2.12837e-13) (5.19193e-14,-3.61739e-14) (-3.94459e-15,-9.74935e-15) (-1.60794e-15,2.75219e-16) (-4.3139e-18,2.23444e-16) (2.84856e-17,5.43874e-18) (1.19051e-18,-3.04394e-18) (-2.87928e-19,-1.69794e-19) (-2.0855e-20,1.99055e-20) (4.8377e-23,1.8692e-21) (4.48883e-23,1.91145e-22) (5.17973e-23,3.14791e-24) (4.42364e-24,-8.14602e-24) (-1.0343e-24,-5.05354e-25) 
  (-3.21411e-29,-1.81268e-30) (2.39107e-30,3.53609e-28) (3.68645e-27,-2.54393e-28) (-4.54829e-27,-3.66836e-26) (-3.45505e-25,6.11628e-26) (6.57908e-25,3.09759e-24) (2.62765e-23,-6.38117e-24) (-4.95052e-23,-2.11195e-22) (-1.62332e-21,3.37282e-22) (1.22364e-21,1.17184e-20) (8.41972e-20,3.66405e-21) (1.72397e-19,-5.60656e-19) (-4.06131e-18,-2.36306e-18) (-2.44123e-17,2.6896e-17) (2.08285e-16,2.21157e-16) (1.60285e-15,-1.43695e-15) (-1.07779e-14,-1.13496e-14) (-5.99665e-14,7.11092e-14) (4.40295e-13,3.26399e-13) (1.12534e-12,-2.47559e-12) (-1.13412e-11,-4.17825e-12) (-4.00358e-12,5.04633e-11) (1.51349e-10,-8.19785e-12) (-1.48363e-10,-4.98602e-10) (-7.03396e-10,5.31047e-10) (9.3528e-10,2.09067e-09) (-9.02419e-12,-2.74783e-09) (1.92938e-09,-5.67796e-09) (8.49016e-09,1.74482e-08) (-3.24465e-08,-2.70395e-08) (2.79522e-08,1.95603e-08) (-2.91386e-08,-1.23063e-08) (2.87176e-08,2.89822e-08) (-2.53081e-08,-6.82953e-09) (5.92675e-08,3.96766e-09) (-1.37575e-10,5.94258e-08) (-3.66056e-08,-1.4288e-08) (4.0804e-08,-3.85125e-08) (1.62622e-08,-1.36941e-08) (-7.32356e-09,-7.27434e-10) (-1.60666e-09,1.17473e-09) (7.0248e-10,1.35465e-09) (-1.47926e-10,2.48259e-10) (-3.67141e-10,-1.09826e-10) (-5.03695e-11,4.16792e-12) (5.24784e-11,-1.48407e-11) (1.00356e-11,-2.26778e-11) (-5.97586e-12,-4.58934e-12) (-1.93492e-12,1.32689e-12) (1.28809e-13,5.36079e-13) (1.14561e-13,1.88556e-15) (6.29899e-15,-2.12055e-14) (-3.20962e-15,-1.88657e-15) (-3.9875e-16,4.24729e-16) (4.6419e-17,6.64227e-17) (9.60892e-18,-4.4181e-18) (-2.79038e-19,-1.19195e-18) (-1.27238e-19,6.26785e-21) (-2.66425e-21,1.13981e-20) (5.85588e-22,6.70927e-22) (7.48194e-23,3.0498e-23) (1.32499e-23,-1.16302e-23) (-8.02931e-25,-3.1054e-24) (-3.88456e-25,8.1081e-26) 
  (-9.78502e-30,5.81795e-30) (7.04739e-29,1.01677e-28) (9.98114e-28,-7.96842e-28) (-8.4648e-27,-9.33749e-27) (-8.23322e-26,8.38382e-26) (7.73086e-25,6.96572e-25) (5.54333e-24,-6.60667e-24) (-5.11614e-23,-4.33231e-23) (-3.23911e-22,3.61257e-22) (2.10711e-21,2.49273e-21) (1.93495e-20,-1.01948e-20) (-1.3576e-20,-1.5735e-19) (-1.3438e-18,-2.48925e-19) (-4.65608e-18,1.09972e-17) (9.36825e-17,4.03904e-17) (3.03728e-16,-6.87995e-16) (-5.15253e-15,-1.69034e-15) (-6.67452e-15,3.13632e-14) (1.8906e-13,1.66681e-14) (-1.08089e-13,-8.99295e-13) (-4.03793e-12,9.32969e-13) (8.20337e-12,1.40926e-11) (4.0577e-11,-3.00818e-11) (-1.34664e-10,-9.46404e-11) (-9.90795e-11,2.47072e-10) (6.99729e-10,3.09021e-10) (-4.58618e-10,-4.98567e-10) (-1.42418e-09,-1.59412e-09) (6.90307e-09,1.26167e-09) (-1.33998e-08,1.81616e-09) (9.74184e-09,-2.10898e-09) (-9.37461e-09,2.98879e-09) (1.264e-08,8.04841e-10) (-8.02256e-09,4.97482e-09) (1.2543e-08,-1.32362e-08) (1.53967e-08,1.22779e-08) (-1.04916e-08,7.28621e-09) (-4.60422e-10,-1.57391e-08) (4.44446e-10,-7.65761e-09) (-1.85069e-09,8.22516e-10) (-1.96e-10,6.8417e-10) (4.5892e-10,1.94745e-10) (5.84722e-11,9.25812e-11) (-9.59145e-11,5.75584e-11) (-1.4513e-11,1.45753e-11) (6.87636e-12,-1.3526e-11) (-2.72045e-12,-7.39348e-12) (-2.40848e-12,1.35133e-13) (-1.87408e-13,7.36953e-13) (1.49023e-13,1.09281e-13) (3.03885e-14,-2.37771e-14) (-2.85224e-15,-6.98224e-15) (-1.27741e-15,1.64775e-16) (-2.09771e-17,2.02069e-16) (2.71945e-17,9.18636e-18) (1.86218e-18,-3.27771e-18) (-3.33079e-19,-2.97864e-19) (-3.80101e-20,2.83393e-20) (1.62512e-21,4.2693e-21) (3.80204e-22,7.01205e-23) (3.02061e-23,-1.5798e-23) (4.05182e-25,-6.04804e-24) (-9.2287e-25,-5.80432e-25) (-8.66303e-26,1.04238e-25) 
  (-1.65294e-30,3.57292e-30) (3.96564e-29,1.47511e-29) (1.19736e-28,-4.1475e-28) (-4.10731e-27,-8.66735e-28) (-5.39461e-27,3.80606e-26) (3.31911e-25,2.79155e-26) (9.9288e-26,-2.6687e-24) (-1.99096e-23,-5.48664e-25) (-6.97444e-24,1.33326e-22) (7.9137e-22,1.86753e-22) (2.74411e-21,-3.96564e-21) (-1.35716e-20,-3.83255e-20) (-4.08841e-19,2.56082e-20) (-2.80233e-19,4.06546e-18) (3.46068e-17,3.04727e-19) (-7.11332e-18,-2.6411e-16) (-1.81812e-15,3.29758e-16) (3.17316e-15,1.05403e-14) (5.70774e-14,-2.89302e-14) (-1.84366e-13,-2.34976e-13) (-9.43209e-13,1.01204e-12) (4.63595e-12,2.21693e-12) (5.39548e-12,-1.56805e-11) (-5.01536e-11,2.46425e-12) (1.23817e-11,8.20167e-11) (2.31756e-10,-7.768e-11) (-1.47824e-10,-3.40293e-11) (-7.56801e-10,1.47293e-10) (1.83986e-09,-1.61477e-09) (-2.39373e-09,3.40442e-09) (1.47863e-09,-2.41075e-09) (-1.63799e-09,2.54395e-09) (3.02045e-09,-2.44029e-09) (-5.93144e-10,3.22406e-09) (-7.38554e-10,-5.38221e-09) (6.17369e-09,-1.38925e-09) (-6.96763e-13,4.05067e-09) (-3.25421e-09,-2.67983e-09) (-1.76468e-09,-1.88462e-09) (-3.86725e-10,4.48492e-10) (8.40438e-11,2.19199e-10) (1.51795e-10,-4.52617e-11) (4.22779e-11,1.14957e-12) (-5.68062e-12,3.08117e-11) (-2.55996e-13,7.55972e-12) (-1.45411e-12,-3.76209e-12) (-2.19842e-12,-1.02928e-12) (-5.424e-13,5.29687e-13) (1.0956e-13,2.1403e-13) (6.02655e-14,-4.55559e-15) (2.81019e-15,-1.24109e-14) (-2.19962e-15,-1.21234e-15) (-3.05835e-16,3.10316e-16) (3.62108e-17,5.90511e-17) (9.44987e-18,-3.07568e-18) (-1.44925e-19,-1.30688e-18) (-1.58094e-19,-1.77171e-20) (-5.57964e-21,1.6307e-20) (1.41701e-21,9.77926e-22) (1.39464e-22,-7.23186e-23) (4.01828e-24,-1.35054e-23) (-1.37549e-24,-1.59936e-24) (-3.58503e-25,7.18303e-26) (-4.52612e-28,4.58153e-26) 
  (2.34388e-31,1.3133e-30) (1.36977e-29,-3.67982e-30) (-4.87085e-29,-1.34538e-28) (-1.24402e-27,5.75529e-28) (6.06659e-27,1.07428e-26) (8.66771e-26,-5.82082e-26) (-4.95522e-25,-6.39043e-25) (-4.36997e-24,3.70174e-24) (2.25187e-23,2.61369e-23) (1.47504e-22,-8.35423e-23) (2.54158e-22,-7.06241e-22) (-4.32138e-21,-1.04979e-20) (-1.32726e-19,3.45638e-20) (3.99816e-19,1.37754e-18) (1.10228e-17,-4.58971e-18) (-4.36628e-17,-8.13291e-17) (-4.8409e-16,3.9013e-16) (2.71126e-15,2.57815e-15) (1.08516e-14,-1.80366e-14) (-9.15148e-14,-3.38926e-14) (-6.62274e-14,4.43937e-13) (1.57737e-12,-2.28392e-13) (-1.5043e-12,-5.10993e-12) (-1.13725e-11,9.52774e-12) (1.70947e-11,2.03937e-11) (3.67271e-11,-6.53397e-11) (-3.47877e-11,1.84851e-12) (-1.03966e-10,2.5749e-10) (-1.98339e-11,-8.20261e-10) (2.50237e-10,1.20787e-09) (-1.82284e-10,-7.59713e-10) (1.00511e-10,9.20591e-10) (1.48648e-10,-1.16253e-09) (6.758e-10,8.66332e-10) (-1.36549e-09,-7.87099e-10) (8.74549e-10,-1.76673e-09) (1.01851e-09,7.25034e-10) (-1.05634e-09,1.88277e-10) (-8.19754e-10,-7.19187e-12) (-5.07454e-11,1.84943e-10) (6.09426e-11,4.07166e-11) (2.70394e-11,-4.05608e-11) (1.01651e-11,-1.20294e-11) (5.3746e-12,6.48506e-12) (1.73654e-12,1.90432e-12) (-9.62711e-13,-3.42466e-13) (-6.81155e-13,2.51169e-13) (-1.67215e-14,2.33318e-13) (6.91714e-14,2.71573e-14) (1.35957e-14,-1.36941e-14) (-1.8477e-15,-3.67438e-15) (-8.05033e-16,1.44861e-16) (-1.57141e-17,1.43331e-16) (2.16058e-17,8.22929e-18) (1.93011e-18,-2.75653e-18) (-3.03476e-19,-3.31162e-19) (-4.82077e-20,2.70995e-20) (1.68642e-21,5.88399e-21) (6.29077e-22,-3.83493e-24) (2.56847e-23,-5.49324e-23) (-2.51389e-24,-5.01843e-24) (-7.36122e-25,-7.12881e-26) (-6.99937e-26,9.91877e-26) (9.68491e-27,1.18647e-26) 
  (3.17184e-31,3.10735e-31) (2.93632e-30,-3.63629e-30) (-3.89843e-29,-2.56437e-29) (-2.03643e-28,3.90978e-28) (3.62877e-27,1.45026e-27) (8.76755e-27,-3.11304e-26) (-2.3939e-25,-4.09336e-26) (-9.78983e-26,1.63002e-24) (8.71921e-24,-5.80855e-25) (-5.01827e-24,-2.73766e-23) (1.63613e-22,-2.02607e-23) (-1.60487e-21,-3.89652e-21) (-4.51282e-20,2.46499e-20) (3.17161e-19,4.03008e-19) (2.84838e-18,-3.04661e-18) (-2.6407e-17,-1.77258e-17) (-7.84189e-17,1.91729e-16) (1.21974e-15,2.80069e-16) (-1.29611e-16,-6.77659e-15) (-3.08637e-14,6.43944e-15) (6.26165e-14,1.27019e-13) (3.64483e-13,-3.25634e-13) (-1.32196e-12,-1.01474e-12) (-1.03295e-12,4.14605e-12) (8.26488e-12,2.48485e-12) (-4.62229e-12,-2.16461e-11) (-1.24411e-11,2.13323e-12) (5.29419e-11,8.27377e-11) (-2.03481e-10,-1.68437e-10) (2.99478e-10,1.8614e-10) (-1.76906e-10,-1.15256e-10) (2.01159e-10,1.98856e-10) (-2.12899e-10,-2.74337e-10) (3.55322e-10,2.00343e-11) (-4.10895e-10,1.76518e-10) (-2.46245e-10,-5.41973e-10) (3.55654e-10,-1.20263e-10) (-1.26039e-10,2.25254e-10) (-1.72155e-10,1.7735e-10) (1.65569e-11,6.37576e-11) (2.22436e-11,2.31535e-13) (-1.53767e-12,-1.43877e-11) (-8.0456e-13,-5.51961e-12) (2.18056e-12,-7.93803e-14) (8.24217e-13,3.43712e-14) (-2.0979e-13,1.28872e-13) (-8.51694e-14,1.92994e-13) (4.36351e-14,5.58023e-14) (2.11167e-14,-7.73419e-15) (3.81809e-16,-6.00728e-15) (-1.19461e-15,-5.21116e-16) (-1.6974e-16,1.98092e-16) (2.49704e-17,3.94767e-17) (7.23109e-18,-2.20812e-18) (-4.33123e-20,-1.11447e-18) (-1.47584e-19,-2.88684e-20) (-7.83649e-21,1.70829e-20) (1.65805e-21,1.3281e-21) (1.81647e-22,-1.30251e-22) (-4.76867e-24,-2.19307e-23) (-1.99375e-24,-8.01739e-25) (-2.06317e-25,1.57155e-25) (5.57417e-27,3.95956e-26) (4.97547e-27,9.19967e-28) 
  (1.43968e-31,2.13228e-32) (6.03186e-32,-1.51778e-30) (-1.49923e-29,1.09462e-30) (2.69579e-29,1.37826e-28) (1.16942e-27,-3.85197e-28) (-4.45591e-27,-8.98621e-27) (-6.03012e-26,4.30192e-26) (3.60006e-25,3.28422e-25) (9.81702e-25,-2.40363e-24) (-1.10352e-23,5.25336e-24) (1.39613e-22,-1.15627e-23) (-1.02607e-21,-1.52556e-21) (-1.32741e-20,1.49498e-20) (1.62431e-19,8.53621e-20) (4.27325e-19,-1.39326e-18) (-1.0721e-17,-9.38967e-19) (8.52819e-18,6.78311e-17) (3.89081e-16,-1.30114e-16) (-1.17517e-15,-1.793e-15) (-7.15103e-15,7.03931e-15) (3.80704e-14,2.11194e-14) (3.76415e-14,-1.43659e-13) (-5.06591e-13,-9.12443e-15) (4.28954e-13,1.13187e-12) (2.63031e-12,-8.8073e-13) (-4.99636e-12,-3.88001e-12) (-4.72099e-12,3.36974e-12) (3.36104e-11,2.86587e-12) (-8.08665e-11,1.21372e-11) (9.43938e-11,-2.37442e-11) (-5.56824e-11,8.25918e-12) (8.571e-11,7.35667e-12) (-1.00337e-10,-1.00628e-11) (7.76117e-11,-8.01193e-11) (-2.7195e-11,1.2174e-10) (-1.6837e-10,-4.49181e-11) (3.29497e-11,-1.04718e-10) (2.29475e-11,5.34218e-11) (2.71582e-12,7.09813e-11) (1.70825e-11,1.46621e-11) (5.80983e-12,-3.45279e-12) (-2.95848e-12,-2.87537e-12) (-1.54093e-12,-1.076e-12) (2.9326e-13,-4.68512e-13) (1.80783e-13,-1.72788e-13) (-4.26613e-15,5.63562e-14) (2.30725e-14,5.4981e-14) (2.07728e-14,3.38757e-15) (3.15547e-15,-5.88193e-15) (-1.12432e-15,-1.45146e-15) (-3.88468e-16,1.14832e-16) (-1.75607e-18,8.15498e-17) (1.40244e-17,4.79801e-18) (1.38975e-18,-1.98647e-18) (-2.31228e-19,-2.78672e-19) (-4.45111e-20,2.13483e-20) (1.25948e-21,6.12346e-21) (7.19926e-22,3.7764e-23) (2.4912e-23,-7.32887e-23) (-6.09093e-24,-5.20968e-24) (-7.51437e-25,2.51121e-25) (-1.69542e-26,8.87382e-26) (1.01356e-26,8.25931e-27) (1.42765e-27,-8.30482e-28) 
  (4.15755e-32,-2.21472e-32) (-2.79742e-31,-4.00524e-31) (-3.54988e-30,3.23763e-30) (3.4388e-29,2.83876e-29) (1.98715e-28,-3.34709e-28) (-2.96647e-27,-1.09135e-27) (-3.08052e-27,2.33562e-26) (1.58414e-25,-2.93947e-26) (-6.3787e-25,-7.93379e-25) (-1.31246e-24,7.42024e-24) (6.58086e-23,-3.78401e-23) (-6.4381e-22,-4.47596e-22) (-2.26938e-21,7.28495e-21) (6.49709e-20,1.96158e-21) (-9.32187e-20,-4.94578e-19) (-3.24826e-18,1.48806e-18) (1.35081e-17,1.77514e-17) (8.36726e-17,-1.01527e-16) (-6.07609e-16,-2.77288e-16) (-6.55093e-16,3.06575e-15) (1.30179e-14,-1.27217e-15) (-1.46191e-14,-4.22259e-14) (-1.21814e-13,8.69575e-14) (2.76633e-13,1.99572e-13) (4.97313e-13,-7.1661e-13) (-1.76504e-12,1.34497e-14) (-7.05195e-13,2.36829e-12) (7.77135e-12,-8.04081e-12) (-1.36257e-11,2.02152e-11) (1.31655e-11,-2.23912e-11) (-1.00458e-11,1.11416e-11) (2.09852e-11,-1.51952e-11) (-2.13005e-11,1.92298e-11) (-3.12917e-12,-3.37302e-11) (2.31869e-11,2.53987e-11) (-4.02013e-11,2.88065e-11) (-1.84891e-11,-2.52493e-11) (1.18902e-11,2.28295e-12) (1.46052e-11,1.29169e-11) (7.40521e-12,2.9615e-13) (1.00192e-12,-1.846e-12) (-1.12129e-12,-9.48087e-14) (-5.93636e-13,1.13115e-13) (-6.67856e-14,-1.25211e-13) (-8.86036e-16,-7.21515e-14) (1.02163e-14,7.30239e-15) (1.54283e-14,5.61657e-15) (5.08117e-15,-3.43602e-15) (-4.5824e-16,-1.89129e-15) (-5.38689e-16,-1.01062e-16) (-6.76137e-17,1.03368e-16) (1.55114e-17,1.96467e-17) (4.32907e-18,-1.58608e-18) (-4.3676e-20,-7.61448e-19) (-1.12472e-19,-2.52177e-20) (-7.32271e-21,1.41104e-20) (1.51699e-21,1.36017e-21) (2.00699e-22,-1.30446e-22) (-7.68592e-24,-2.50214e-23) (-2.76978e-24,-1.66399e-25) (-1.4902e-25,2.39617e-25) (1.56568e-26,2.68591e-26) (4.23618e-27,-2.29476e-28) (1.72908e-28,-5.03767e-28) 
  (6.39903e-33,-1.36743e-32) (-1.48873e-31,-4.66409e-32) (-2.3742e-31,1.51137e-30) (1.41888e-29,-1.03369e-31) (-2.3671e-29,-1.2211e-28) (-9.36324e-28,4.10411e-28) (4.998e-27,6.11018e-27) (2.88001e-26,-5.08009e-26) (-4.33012e-25,-1.29712e-26) (1.81617e-24,3.14923e-24) (1.71617e-23,-2.90551e-23) (-3.10454e-22,-4.61138e-23) (4.82685e-22,2.76763e-21) (2.03564e-20,-9.90053e-21) (-1.09164e-19,-1.30895e-19) (-6.70354e-19,9.51966e-19) (6.65729e-18,2.67196e-18) (5.08075e-18,-4.09584e-17) (-2.03291e-16,2.81792e-17) (3.56663e-16,8.90306e-16) (2.95318e-15,-2.47509e-15) (-1.06429e-14,-7.94425e-15) (-1.34056e-14,4.08766e-14) (9.65114e-14,5.64289e-15) (-1.33244e-14,-2.66515e-13) (-3.92777e-13,2.89782e-13) (4.18409e-13,8.60629e-13) (-3.4504e-13,-3.55529e-12) (1.56954e-12,6.83227e-12) (-1.6528e-12,-6.50352e-12) (-2.92087e-13,4.04925e-12) (1.60501e-12,-7.51114e-12) (1.62408e-13,8.0119e-12) (-8.16441e-12,-5.7377e-12) (9.32495e-12,-1.30463e-12) (-9.01666e-13,1.35822e-11) (-8.70895e-12,-3.2316e-14) (1.42001e-12,-1.83805e-12) (5.0955e-12,-4.26894e-13) (1.82599e-12,-1.44503e-12) (-4.06455e-14,-6.6682e-13) (-2.43404e-13,1.62112e-13) (-1.04556e-13,1.5382e-13) (-3.89403e-14,8.74126e-16) (-1.49664e-14,-1.30949e-14) (2.48036e-15,-1.39545e-15) (3.89964e-15,-2.0654e-15) (3.6392e-16,-1.71507e-15) (-4.60707e-16,-3.14767e-16) (-1.37148e-16,8.29937e-17) (4.79809e-18,3.66443e-17) (7.38103e-18,1.56867e-18) (7.17685e-19,-1.20994e-18) (-1.56883e-19,-1.75691e-19) (-3.25591e-20,1.5357e-20) (8.52961e-22,4.95152e-21) (6.48593e-22,5.85731e-23) (2.74592e-23,-7.28168e-23) (-6.92789e-24,-5.18773e-24) (-7.78243e-25,5.17322e-25) (1.22814e-26,9.66052e-26) (9.93299e-27,3.49538e-27) (9.68582e-28,-9.6123e-28) (-6.35137e-29,-1.57326e-28) 
  (-1.00669e-33,-4.69611e-33) (-4.64274e-32,1.74372e-32) (2.43818e-31,4.21408e-31) (3.44847e-30,-2.95242e-30) (-3.20023e-29,-2.44636e-29) (-1.32976e-28,3.11954e-28) (2.72948e-27,2.81393e-28) (-5.86253e-27,-2.10236e-26) (-1.34666e-25,1.14368e-25) (1.39528e-24,6.14534e-25) (-1.04433e-25,-1.34878e-23) (-1.10838e-22,4.15969e-23) (6.25721e-22,7.75789e-22) (4.42583e-21,-6.32091e-21) (-5.30212e-20,-1.92208e-20) (-2.83716e-20,3.71596e-19) (2.23453e-18,-3.82494e-19) (-5.48282e-18,-1.14341e-17) (-4.72181e-17,4.04911e-17) (2.38128e-16,1.60219e-16) (3.05294e-16,-1.07404e-15) (-3.88368e-15,-1.47049e-16) (3.66027e-15,1.15008e-14) (2.43048e-14,-1.33495e-14) (-5.18937e-14,-6.00286e-14) (-4.63561e-14,1.28614e-13) (3.23448e-13,1.15877e-13) (-8.90904e-13,-6.44522e-13) (1.67509e-12,9.92697e-13) (-1.42664e-12,-8.89897e-13) (6.1713e-13,9.44212e-13) (-1.15516e-12,-1.90774e-12) (1.72112e-12,1.37266e-12) (-2.76106e-12,7.2428e-13) (1.13398e-12,-2.30324e-12) (2.65322e-12,2.48387e-12) (-1.41599e-12,1.89878e-12) (-2.935e-13,-3.47031e-13) (8.05478e-13,-9.94244e-13) (1.15425e-13,-6.88367e-13) (-1.3083e-13,-1.68972e-13) (-2.41187e-14,6.80506e-14) (9.81186e-15,5.40312e-14) (-5.16183e-15,1.04818e-14) (-5.19704e-15,7.67795e-16) (-1.03909e-16,-7.07444e-16) (2.70538e-16,-1.12828e-15) (-2.64762e-16,-4.14178e-16) (-1.55986e-16,2.17927e-17) (-1.33205e-17,4.40154e-17) (8.11705e-18,7.20539e-18) (1.97586e-18,-1.04686e-18) (-6.3844e-20,-4.16548e-19) (-7.04534e-20,-1.18358e-20) (-4.95228e-21,9.86644e-21) (1.14442e-21,1.05908e-21) (1.73679e-22,-1.07591e-22) (-6.79842e-24,-2.38449e-23) (-2.80151e-24,-2.41647e-26) (-1.01749e-25,2.89645e-25) (2.34886e-26,2.26898e-26) (3.28179e-27,-1.22382e-27) (3.13554e-29,-4.33443e-28) (-4.74941e-29,-2.4361e-29) 
  (-1.154e-33,-9.87975e-34) (-8.17254e-33,1.34281e-32) (1.44765e-31,5.55105e-32) (2.40941e-31,-1.44043e-30) (-1.31567e-29,8.28929e-31) (3.67429e-29,1.08098e-28) (7.76337e-28,-5.7138e-28) (-6.73435e-27,-4.41336e-27) (-1.3332e-26,6.65731e-26) (5.75421e-25,-1.12395e-25) (-2.67973e-24,-4.25646e-24) (-2.6681e-23,3.30522e-23) (3.19176e-22,1.22161e-22) (2.15033e-22,-2.55958e-21) (-1.78766e-20,3.51521e-21) (5.31107e-20,1.04481e-19) (5.22896e-19,-4.69328e-19) (-3.25856e-18,-1.99729e-18) (-5.21253e-18,1.78276e-17) (8.40215e-17,-7.04469e-19) (-9.93054e-17,-3.03231e-16) (-9.39541e-16,6.0362e-16) (2.64282e-15,2.01109e-15) (3.86601e-15,-7.04907e-15) (-2.25428e-14,-4.48726e-15) (8.69894e-15,3.86167e-14) (1.04868e-13,-4.98681e-14) (-3.19541e-13,6.7352e-14) (5.04614e-13,-1.37715e-13) (-4.03051e-13,7.56006e-14) (3.04006e-13,1.04164e-13) (-6.12441e-13,-1.57119e-13) (5.82202e-13,-1.31293e-13) (-3.39272e-13,7.1749e-13) (-3.43343e-13,-6.06764e-13) (9.33072e-13,-1.27559e-13) (1.81332e-13,6.03439e-13) (-9.96264e-14,7.54983e-14) (-3.72914e-14,-3.02191e-13) (-1.10584e-13,-1.66592e-13) (-6.49304e-14,-1.80791e-14) (4.1671e-15,1.64543e-14) (1.26629e-14,9.07212e-15) (1.97589e-15,3.11117e-15) (-6.68844e-16,1.15906e-15) (-1.94799e-16,-5.17422e-17) (-1.75112e-16,-2.42658e-16) (-1.32171e-16,-2.86857e-17) (-2.78299e-17,3.38255e-17) (5.53876e-18,1.17099e-17) (3.1298e-18,2.00564e-20) (2.43583e-19,-6.04473e-19) (-9.25783e-20,-8.25404e-20) (-1.85527e-20,1.04451e-20) (6.71404e-22,3.25782e-21) (4.73497e-22,4.23044e-23) (2.26318e-23,-5.87449e-23) (-6.16541e-24,-4.69325e-24) (-7.1842e-25,5.23107e-25) (2.99464e-26,9.39302e-26) (1.06189e-26,1.0307e-27) (5.73564e-28,-9.88441e-28) (-8.11779e-29,-1.10186e-28) (-1.6121e-29,3.8827e-30) 
  (-4.77407e-34,-2.69952e-35) (5.76506e-34,4.93577e-33) (4.70376e-32,-1.50141e-32) (-2.34678e-31,-4.08435e-31) (-3.13681e-30,2.98585e-30) (3.30012e-29,1.98342e-29) (7.97158e-29,-3.25867e-28) (-2.87178e-27,2.66056e-28) (1.04942e-26,2.24202e-26) (1.49537e-25,-1.50556e-25) (-1.60698e-24,-7.69762e-25) (-1.90515e-24,1.44898e-23) (1.11917e-22,-1.98268e-23) (-3.69414e-22,-7.47884e-22) (-4.2211e-21,3.90424e-21) (3.09602e-20,1.87774e-20) (5.67007e-20,-2.05694e-19) (-1.13137e-18,3.01141e-20) (1.60998e-18,5.21362e-18) (1.97491e-17,-1.37944e-17) (-7.10115e-17,-5.537e-17) (-1.1906e-16,2.91164e-16) (9.00622e-16,4.80934e-17) (-1.85622e-16,-2.33209e-15) (-5.84356e-15,2.87898e-15) (8.50651e-15,8.32506e-15) (1.22202e-14,-3.52557e-14) (-4.81925e-14,8.03447e-14) (6.6649e-14,-1.18611e-13) (-6.07433e-14,7.68432e-14) (8.6814e-14,-3.24993e-14) (-1.49631e-13,9.02488e-14) (6.82369e-14,-1.44881e-13) (9.03877e-14,1.9474e-13) (-1.87348e-13,-1.69917e-14) (1.22009e-13,-2.03121e-13) (1.54231e-13,5.57988e-14) (1.51523e-14,4.12594e-14) (-5.45076e-14,-4.13774e-14) (-5.35178e-14,-1.20382e-14) (-1.90156e-14,8.14773e-15) (2.63788e-15,2.86101e-15) (4.20588e-15,-5.97882e-16) (1.16087e-15,6.32026e-17) (1.37059e-16,3.03266e-16) (-4.04674e-17,4.25727e-17) (-7.57179e-17,-5.61884e-18) (-3.04724e-17,2.01616e-17) (7.33864e-19,1.19867e-17) (3.31698e-18,1.36496e-18) (6.67831e-19,-5.83125e-19) (-5.90746e-20,-1.77319e-19) (-3.5873e-20,-1.23764e-21) (-2.28567e-21,5.80377e-21) (7.56405e-22,6.31418e-22) (1.1975e-22,-7.71547e-23) (-5.3496e-24,-1.8299e-23) (-2.37688e-24,-1.07127e-26) (-8.16534e-26,2.6415e-25) (2.53198e-26,1.78909e-26) (2.86289e-27,-1.83857e-27) (-5.70654e-29,-3.61115e-28) (-4.13854e-29,-1.00127e-29) (-2.9889e-30,4.11447e-30) 
  (-1.24239e-34,8.36158e-35) (1.0944e-33,1.11909e-33) (8.79806e-33,-1.29901e-32) (-1.41078e-31,-5.56022e-32) (-1.86936e-31,1.40512e-30) (1.27534e-29,-1.72076e-30) (-4.71921e-29,-1.04297e-28) (-7.41492e-28,6.70763e-28) (7.50984e-27,4.26425e-27) (1.40189e-26,-7.19823e-26) (-6.01391e-25,7.32711e-26) (2.0126e-24,4.41425e-24) (2.74723e-23,-2.44378e-23) (-2.24271e-22,-1.39804e-22) (-4.63638e-22,1.71337e-21) (1.09821e-20,-2.01969e-22) (-1.92197e-20,-6.05004e-20) (-2.70982e-19,1.87712e-19) (1.22302e-18,9.92332e-19) (2.39237e-18,-6.33798e-18) (-2.50432e-17,-1.7596e-18) (1.91723e-17,8.47052e-17) (2.10186e-16,-1.2292e-16) (-4.24285e-16,-5.28139e-16) (-8.22175e-16,1.62085e-15) (3.60888e-15,6.17943e-16) (-5.10399e-15,-1.02779e-14) (7.00724e-15,2.50407e-14) (-9.16868e-15,-3.30569e-14) (3.7808e-16,2.31571e-14) (1.26073e-14,-2.34912e-14) (-1.01323e-14,4.59583e-14) (-1.95893e-14,-3.78488e-14) (5.47167e-14,1.43114e-14) (-3.25987e-14,3.82305e-14) (-2.04732e-14,-5.41952e-14) (3.4857e-14,-2.30309e-14) (1.47565e-14,2.32139e-15) (-1.42055e-14,1.99664e-15) (-1.23029e-14,7.54203e-15) (-2.73658e-15,5.49732e-15) (8.47218e-16,4.04553e-16) (6.94968e-16,-8.70356e-16) (2.37866e-16,-2.65904e-16) (8.19511e-17,1.17975e-17) (3.89282e-18,1.60969e-17) (-1.31475e-17,1.37228e-17) (-1.72527e-18,9.54561e-18) (2.36832e-18,2.22134e-18) (9.17703e-19,-3.36222e-19) (3.06483e-20,-2.44912e-19) (-4.52471e-20,-2.71371e-20) (-8.06038e-21,6.28528e-21) (5.50358e-22,1.71103e-21) (2.87034e-22,5.76746e-24) (1.37312e-23,-3.96693e-23) (-4.58565e-24,-3.34744e-24) (-5.72328e-25,4.30701e-25) (2.85772e-26,7.94492e-26) (9.55495e-27,-3.1397e-28) (3.48993e-28,-1.00224e-27) (-8.50117e-29,-7.69766e-29) (-1.17536e-29,5.73123e-30) (1.12532e-31,1.53537e-30) 
  (-1.53027e-35,4.40417e-35) (4.85173e-34,7.13428e-35) (-2.99625e-34,-4.94984e-33) (-4.65532e-32,1.35759e-32) (2.30864e-31,3.97273e-31) (2.98928e-30,-3.00007e-30) (-3.34045e-29,-1.84273e-29) (-7.04976e-29,3.28434e-28) (2.89085e-27,-2.5762e-28) (-9.37096e-27,-2.25432e-26) (-1.53008e-25,1.27198e-25) (1.30788e-24,8.52483e-25) (3.24401e-24,-1.11318e-23) (-8.17419e-23,5.0621e-25) (1.59675e-22,5.12346e-22) (2.7184e-21,-1.81741e-21) (-1.43703e-20,-1.16744e-20) (-3.52971e-20,8.76558e-20) (4.44553e-19,3.91199e-20) (-4.39381e-19,-1.8199e-18) (-5.98787e-18,3.45107e-18) (1.73487e-17,1.58988e-17) (2.97878e-17,-5.86461e-17) (-1.86259e-16,-5.40859e-17) (8.16339e-17,4.96029e-16) (1.00374e-15,-5.13977e-16) (-3.22522e-15,-1.0549e-15) (6.1566e-15,3.31118e-15) (-7.24695e-15,-4.23896e-15) (3.42195e-15,4.31294e-15) (-1.92184e-15,-7.3066e-15) (7.08187e-15,1.0129e-14) (-1.10875e-14,-1.92121e-15) (1.17407e-14,-8.54917e-15) (3.11625e-15,1.28547e-14) (-1.31797e-14,-4.02778e-15) (5.84675e-16,-1.03952e-14) (3.22016e-15,-3.39308e-15) (-1.68493e-15,2.15538e-15) (-8.82098e-16,3.53357e-15) (4.5701e-16,1.69855e-15) (2.6107e-16,2.80668e-17) (-2.05223e-17,-2.79747e-16) (-1.34525e-17,-1.04631e-16) (1.31579e-17,-1.6797e-17) (4.1018e-18,1.59694e-18) (5.77386e-19,4.66673e-18) (1.50658e-18,2.03607e-18) (8.66021e-19,-8.56554e-21) (1.19953e-19,-2.33299e-19) (-3.86011e-20,-5.54617e-20) (-1.44458e-20,2.52644e-21) (-5.93282e-22,2.80374e-21) (4.29111e-22,2.74943e-22) (6.50892e-23,-5.04007e-23) (-4.0082e-24,-1.14923e-23) (-1.66272e-24,4.79785e-26) (-5.71535e-26,2.04361e-25) (2.12248e-26,1.38201e-26) (2.24644e-27,-1.82452e-27) (-1.04371e-28,-3.0703e-28) (-3.52224e-29,-2.14909e-30) (-1.65921e-30,3.59775e-30) (3.20029e-31,3.30379e-31) 
  (4.30175e-36,1.37529e-35) (1.34125e-34,-7.25409e-35) (-1.00708e-33,-1.18396e-33) (-9.18926e-33,1.22896e-32) (1.35167e-31,5.75147e-32) (2.01658e-31,-1.3528e-30) (-1.23161e-29,1.49921e-30) (4.26988e-29,1.0096e-28) (7.3013e-28,-5.98976e-28) (-6.53272e-27,-4.39497e-27) (-1.8831e-26,6.05381e-26) (4.88735e-25,3.56051e-27) (-9.98943e-25,-3.42735e-24) (-2.07154e-23,1.34709e-23) (1.21972e-22,1.02111e-22) (3.75779e-22,-8.78051e-22) (-5.27307e-21,-5.20038e-22) (5.36108e-21,2.61172e-20) (1.08402e-19,-6.04341e-20) (-3.76532e-19,-3.4308e-19) (-8.23536e-19,1.68686e-18) (6.21092e-18,8.93156e-19) (-1.733e-18,-1.77675e-17) (-5.16006e-17,1.81825e-17) (9.83595e-17,9.78814e-17) (1.39799e-16,-3.12198e-16) (-8.60637e-16,4.43259e-16) (1.73969e-15,-5.43582e-16) (-1.94625e-15,4.51374e-16) (1.29071e-15,3.52002e-16) (-1.79823e-15,-1.07483e-15) (3.14678e-15,3.73721e-16) (-2.1556e-15,2.00575e-15) (1.84316e-16,-3.63474e-15) (3.15045e-15,1.33151e-15) (-2.58141e-15,1.88438e-15) (-1.94782e-15,-1.62641e-15) (-2.2403e-16,-1.34627e-15) (2.10538e-17,4.4885e-16) (4.48887e-16,7.58392e-16) (4.09743e-16,2.61484e-16) (7.8502e-17,-2.62293e-17) (-4.8994e-17,-4.67896e-17) (-2.45732e-17,-1.72091e-17) (-2.23322e-18,-5.38719e-18) (9.09569e-19,-6.09098e-19) (9.76156e-19,6.09707e-19) (6.47052e-19,7.18905e-20) (1.61982e-19,-1.60338e-19) (-1.87256e-20,-6.68492e-20) (-1.77383e-20,-4.08808e-21) (-2.52395e-21,3.12201e-21) (3.75885e-22,6.96669e-22) (1.41195e-22,-1.74855e-23) (5.28626e-24,-2.26311e-23) (-2.93782e-24,-1.85369e-24) (-3.69419e-25,3.06011e-25) (2.31393e-26,5.73506e-26) (7.4478e-27,-5.54255e-28) (2.02814e-28,-8.36616e-28) (-8.12148e-29,-5.34203e-29) (-8.72637e-30,6.11639e-30) (2.90624e-31,1.14755e-30) (1.34816e-31,1.48946e-32) 
  (3.5475e-36,2.62687e-36) (2.01061e-35,-4.24414e-35) (-4.68932e-34,-1.1109e-34) (-4.69709e-35,4.79188e-33) (4.50299e-32,-1.03554e-32) (-1.97678e-31,-3.85139e-31) (-2.92418e-30,2.64067e-30) (2.93684e-29,1.87206e-29) (8.54865e-29,-2.86177e-28) (-2.46948e-27,-2.03666e-29) (5.37154e-27,1.89128e-26) (1.25906e-25,-8.01612e-26) (-8.11831e-25,-7.03959e-25) (-2.97208e-24,6.6773e-24) (4.59255e-23,5.56982e-24) (-4.83516e-23,-2.69374e-22) (-1.31571e-21,6.97965e-22) (5.2621e-21,5.20682e-21) (1.52003e-20,-3.02877e-20) (-1.35195e-19,-2.00101e-20) (6.98747e-20,4.97858e-19) (1.49092e-18,-7.14423e-19) (-3.01224e-18,-3.82472e-18) (-8.63801e-18,1.25008e-17) (3.78944e-17,6.10496e-18) (-2.81261e-17,-9.72906e-17) (-8.05525e-17,2.54698e-16) (2.13e-16,-4.093e-16) (-2.62684e-16,3.81913e-16) (3.12872e-16,-1.20426e-16) (-5.48027e-16,1.43779e-16) (5.87505e-16,-5.35161e-16) (7.28021e-17,7.58253e-16) (-6.6735e-16,-5.90441e-16) (7.50124e-16,-4.33402e-16) (3.33061e-18,7.24921e-16) (-5.87649e-16,1.42161e-16) (-3.29223e-16,-1.81246e-16) (2.78073e-17,4.83491e-17) (1.9737e-16,5.17685e-17) (1.2748e-16,-2.36219e-17) (1.7074e-17,-2.03172e-17) (-1.56383e-17,-6.98848e-19) (-8.04292e-18,1.65449e-18) (-1.65086e-18,-2.59675e-19) (-4.14963e-21,-2.55127e-19) (2.63387e-19,-8.99798e-20) (1.24101e-19,-1.08503e-19) (7.73711e-22,-5.91827e-20) (-1.54915e-20,-9.41467e-21) (-4.20647e-21,2.37072e-21) (4.5749e-23,1.08175e-21) (2.00997e-22,7.77861e-23) (2.67079e-23,-2.85913e-23) (-2.84784e-24,-5.80103e-24) (-9.70187e-25,1.09981e-25) (-2.87435e-26,1.3316e-25) (1.53247e-26,8.9368e-27) (1.61603e-27,-1.44246e-27) (-1.01479e-28,-2.30464e-28) (-2.85333e-29,2.24594e-30) (-9.01484e-31,3.02915e-30) (2.7838e-31,2.10038e-31) (3.30981e-32,-2.15183e-32) 
  (1.33813e-36,1.96485e-38) (-2.57765e-36,-1.40671e-35) (-1.36397e-34,5.61685e-35) (8.46357e-34,1.20718e-33) (9.49777e-33,-1.06671e-32) (-1.18799e-31,-6.25573e-32) (-2.80632e-31,1.19051e-30) (1.0791e-29,-3.23171e-31) (-2.72189e-29,-8.79633e-29) (-6.33653e-28,4.11233e-28) (4.49687e-27,3.89424e-27) (1.84287e-26,-4.05656e-26) (-3.13552e-25,-4.321e-26) (3.38503e-25,2.09061e-24) (1.18365e-23,-5.85913e-24) (-5.31971e-23,-5.56124e-23) (-1.95684e-22,3.62048e-22) (1.98588e-21,3.80853e-22) (-1.18828e-21,-9.01436e-21) (-3.27171e-20,1.54934e-20) (8.86686e-20,9.88259e-20) (2.23739e-19,-3.70101e-19) (-1.26029e-18,-4.25416e-19) (1.06889e-19,4.15867e-18) (9.48958e-18,-4.81435e-18) (-2.4568e-17,-1.56911e-17) (3.29368e-17,6.33979e-17) (-3.35216e-17,-1.08477e-16) (1.23806e-17,1.0457e-16) (4.49254e-17,-7.35469e-17) (-7.18589e-17,1.30862e-16) (-7.60619e-18,-1.95223e-16) (1.64243e-16,1.03792e-16) (-2.10007e-16,3.82279e-17) (2.79062e-17,-2.12719e-16) (1.33371e-16,9.13341e-17) (-5.44046e-17,1.29849e-16) (-9.1229e-17,3.73291e-17) (-2.85849e-19,9.29021e-18) (3.90343e-17,-2.24335e-17) (1.96226e-17,-2.70285e-17) (5.42022e-19,-8.19433e-18) (-2.75597e-18,2.07659e-18) (-1.16475e-18,1.82615e-18) (-3.34633e-19,3.52199e-19) (-5.07011e-20,-2.59808e-20) (2.33396e-20,-6.20617e-20) (7.70496e-22,-4.11298e-20) (-1.05707e-20,-1.08788e-20) (-4.57193e-21,9.71134e-22) (-3.90494e-22,1.20007e-21) (2.00025e-22,2.06858e-22) (5.45291e-23,-1.93555e-23) (5.51018e-25,-1.05898e-23) (-1.61294e-24,-7.30562e-25) (-1.89936e-25,1.92462e-25) (1.68239e-26,3.41976e-26) (4.96649e-27,-6.72121e-28) (1.13619e-28,-6.07847e-28) (-6.35642e-29,-3.48459e-29) (-6.12761e-30,5.57775e-30) (3.41101e-31,8.55704e-31) (1.01239e-31,-2.74677e-33) (3.4834e-33,-1.07947e-32) 
  (3.30867e-37,-2.26667e-37) (-3.07477e-36,-3.00671e-36) (-2.38671e-35,3.75821e-35) (4.19793e-34,1.51936e-34) (5.1479e-34,-4.30624e-33) (-4.05282e-32,4.86087e-33) (1.33378e-31,3.46866e-31) (2.65575e-30,-1.90936e-30) (-2.15238e-29,-1.74903e-29) (-9.02003e-29,2.07003e-28) (1.74429e-27,2.31033e-28) (-1.99386e-27,-1.2867e-26) (-8.24694e-26,3.92361e-26) (4.07045e-25,4.43284e-25) (1.86349e-24,-3.19954e-24) (-2.07374e-23,-4.62721e-24) (1.0405e-23,1.11383e-22) (4.9982e-22,-2.12916e-22) (-1.59165e-21,-1.79626e-21) (-4.88705e-21,8.11695e-21) (3.35265e-20,8.60557e-21) (-3.26477e-21,-1.12801e-19) (-3.49945e-19,9.44595e-20) (6.87715e-19,8.90505e-19) (1.30782e-18,-2.64034e-18) (-8.03778e-18,1.34186e-18) (1.76646e-17,5.66092e-18) (-2.38491e-17,-1.3056e-17) (1.71645e-17,1.6167e-17) (-3.13686e-18,-2.21753e-17) (1.22026e-17,3.63443e-17) (-3.7636e-17,-2.8488e-17) (4.59054e-17,-1.63374e-17) (-2.30679e-17,4.44942e-17) (-3.65169e-17,-3.68568e-17) (3.30435e-17,-1.35046e-17) (1.66362e-17,2.7386e-17) (-7.22551e-18,2.36968e-17) (5.15637e-19,4.86285e-18) (2.56537e-18,-9.04064e-18) (-1.14257e-18,-8.23535e-18) (-1.40242e-18,-1.97599e-18) (-2.00225e-19,6.96879e-19) (1.20971e-19,5.37772e-19) (2.17564e-20,1.37731e-19) (-9.79986e-21,8.82807e-21) (-7.61156e-21,-1.34867e-20) (-7.38393e-21,-6.91886e-21) (-3.83639e-21,-3.63675e-23) (-6.74284e-22,9.81131e-22) (1.36022e-22,2.95411e-22) (7.51908e-23,5.41004e-24) (7.55704e-24,-1.33308e-23) (-1.71622e-24,-2.25528e-24) (-4.61301e-25,1.26225e-25) (-7.10178e-27,7.34691e-26) (9.50542e-27,4.48071e-27) (9.71924e-28,-1.00081e-27) (-7.95536e-29,-1.54573e-28) (-2.03003e-29,3.1754e-30) (-4.05148e-31,2.32581e-30) (2.28621e-31,1.32168e-31) (2.2206e-32,-1.86455e-32) (-1.1523e-33,-3.00425e-33) 
  (4.20106e-38,-1.11015e-37) (-1.25826e-36,-2.11176e-37) (5.41061e-37,1.32281e-35) (1.28633e-34,-3.38362e-35) (-6.00307e-34,-1.14593e-33) (-9.17224e-33,8.00265e-33) (9.0701e-32,6.33451e-32) (3.38961e-31,-9.08932e-31) (-8.13875e-30,-7.78336e-31) (1.14183e-29,6.50687e-29) (4.58469e-28,-2.22424e-28) (-2.5043e-27,-2.76346e-27) (-1.33478e-26,2.21208e-26) (1.62922e-25,4.04473e-26) (-6.02295e-26,-1.01789e-24) (-5.37309e-24,2.08391e-24) (1.8878e-23,2.32224e-23) (7.81427e-23,-1.20456e-22) (-6.03912e-22,-1.57356e-22) (1.02838e-22,2.44976e-21) (8.43799e-21,-2.90844e-21) (-1.65935e-20,-2.43577e-20) (-6.36981e-20,7.462e-20) (2.89617e-19,8.31548e-20) (-1.58688e-19,-7.94859e-19) (-1.36201e-18,1.74392e-18) (4.18096e-18,-2.10774e-18) (-6.13377e-18,1.62413e-18) (5.23688e-18,4.27332e-19) (-4.41238e-18,-3.75823e-18) (8.81256e-18,3.81582e-18) (-1.08941e-17,2.75447e-18) (3.87167e-18,-1.13464e-17) (4.95154e-18,1.04419e-17) (-1.21591e-17,1.44278e-18) (1.35784e-18,-7.76017e-18) (7.1145e-18,5.22531e-19) (3.32776e-18,4.98025e-18) (1.30708e-18,1.3695e-18) (-8.51833e-19,-1.62119e-18) (-1.5767e-18,-1.2303e-18) (-6.62926e-19,-1.61891e-19) (4.18958e-20,1.40528e-19) (1.13979e-19,7.31333e-20) (3.34928e-20,1.99093e-20) (1.48637e-21,3.25432e-21) (-3.45872e-21,-6.77599e-22) (-2.44392e-21,2.08876e-22) (-6.76533e-22,6.77785e-22) (4.81523e-23,2.95776e-22) (7.64746e-23,3.14538e-23) (1.53568e-23,-1.19766e-23) (-8.03359e-25,-3.92299e-24) (-7.30045e-25,-1.5921e-25) (-7.2786e-26,1.04549e-25) (1.10419e-26,1.65163e-26) (2.77771e-27,-6.67566e-28) (3.9053e-29,-3.80813e-28) (-4.37185e-29,-2.01902e-29) (-3.9399e-30,4.17156e-30) (3.10472e-31,5.85241e-31) (7.37584e-32,-1.05603e-32) (1.64687e-33,-8.0175e-33) (-7.77981e-34,-4.55151e-34) 
  (-8.25188e-39,-3.36746e-38) (-3.38453e-37,1.57323e-37) (2.31902e-36,3.10788e-36) (2.55694e-35,-2.94309e-35) (-3.34169e-34,-1.792e-34) (-9.15963e-34,3.44352e-33) (3.22964e-32,6.11301e-34) (-6.46993e-32,-2.74475e-31) (-2.08322e-30,1.11362e-30) (1.30336e-29,1.37446e-29) (7.37123e-29,-1.24498e-28) (-1.01529e-27,-2.59309e-28) (3.08092e-28,7.16516e-27) (4.33129e-26,-1.54768e-26) (-1.66459e-25,-2.20055e-25) (-8.81164e-25,1.25902e-24) (7.53395e-24,2.31782e-24) (-6.09522e-25,-3.73368e-23) (-1.5136e-22,5.21945e-23) (3.66278e-22,5.09941e-22) (1.4022e-21,-1.8014e-21) (-7.09773e-21,-3.02051e-21) (-2.51641e-21,2.61814e-20) (7.49851e-20,-2.79765e-20) (-1.68416e-19,-1.42046e-19) (4.94057e-20,5.82004e-19) (3.74756e-19,-1.08767e-18) (-7.73056e-19,1.22163e-18) (9.89642e-19,-6.3921e-19) (-1.47661e-18,7.58321e-20) (2.12509e-18,-1.00176e-18) (-1.07219e-18,2.41493e-18) (-1.55175e-18,-2.43727e-18) (2.57161e-18,5.16019e-19) (-1.46249e-18,2.40984e-18) (-1.31797e-18,-1.15516e-18) (9.78757e-19,-1.20997e-18) (1.39023e-18,1.32709e-19) (6.0431e-19,3.13203e-20) (-3.04588e-19,-1.13029e-19) (-4.61785e-19,5.13605e-20) (-1.62094e-19,8.73148e-20) (2.02506e-20,2.19595e-20) (3.14947e-20,-6.34e-21) (1.00303e-20,-3.25137e-21) (1.11658e-21,-2.68017e-23) (-6.12964e-22,4.75134e-22) (-3.53046e-22,4.67105e-22) (3.80078e-24,2.35849e-22) (5.97307e-23,4.46318e-23) (1.94125e-23,-7.34628e-24) (8.42878e-25,-4.89083e-24) (-8.23852e-25,-6.22901e-25) (-1.71188e-25,9.21891e-26) (3.02397e-27,3.3339e-26) (5.05064e-27,1.52176e-27) (4.66871e-28,-6.07295e-28) (-5.58453e-29,-8.72482e-29) (-1.27949e-29,3.03514e-30) (-1.51128e-31,1.57223e-30) (1.67144e-31,7.50728e-32) (1.43082e-32,-1.49686e-32) (-1.02371e-33,-2.0354e-33) (-2.4682e-34,3.55957e-35) 
  (-7.41791e-39,-6.69268e-39) (-5.53297e-38,9.23172e-38) (1.05639e-36,3.67828e-37) (1.36937e-36,-1.1161e-35) (-1.08722e-34,1.08435e-35) (3.31915e-34,9.69368e-34) (7.79837e-33,-4.99114e-33) (-5.8726e-32,-5.49671e-32) (-3.17526e-31,5.89557e-31) (5.19223e-30,1.19564e-30) (-2.05328e-30,-4.02636e-29) (-2.72887e-28,9.53241e-29) (1.15235e-27,1.57927e-27) (7.3936e-27,-9.93776e-27) (-6.93512e-26,-2.40208e-26) (-8.26509e-27,4.03049e-25) (1.95852e-24,-5.86745e-25) (-5.44771e-24,-7.86017e-24) (-2.47571e-23,3.21607e-23) (1.48444e-22,5.76424e-23) (5.17216e-23,-5.78735e-22) (-1.9904e-21,3.49885e-22) (3.48695e-21,6.03916e-21) (1.14155e-20,-1.77411e-20) (-5.89148e-20,-7.52559e-22) (1.11267e-19,1.00641e-19) (-1.15961e-19,-2.49858e-19) (5.45104e-20,3.17733e-19) (9.22313e-20,-2.51878e-19) (-2.48238e-19,2.74064e-19) (1.50585e-19,-5.41644e-19) (2.91934e-19,5.41117e-19) (-6.7717e-19,-7.53395e-20) (4.33543e-19,-3.96269e-19) (2.24809e-19,5.91769e-19) (-3.76095e-19,1.19958e-19) (-9.85778e-20,-3.18954e-19) (2.20036e-19,-2.24667e-19) (1.2803e-19,-1.16727e-19) (-4.7604e-20,1.46114e-20) (-6.58791e-20,8.06506e-20) (-1.548e-20,4.5179e-20) (6.03935e-21,3.08483e-21) (4.2385e-21,-6.01247e-21) (1.14532e-21,-2.5113e-21) (1.75887e-22,-3.092e-22) (-1.13072e-23,1.62911e-22) (2.59889e-23,1.35016e-22) (4.19378e-23,3.9075e-23) (1.81859e-23,-2.38033e-24) (2.25778e-24,-4.62441e-24) (-6.7402e-25,-1.05043e-24) (-2.622e-25,2.04198e-26) (-1.78278e-26,4.66634e-26) (6.18005e-27,6.09787e-27) (1.27327e-27,-5.37286e-28) (-5.52151e-30,-2.02584e-28) (-2.61906e-29,-8.88039e-30) (-2.1983e-30,2.77671e-30) (2.30455e-31,3.61552e-31) (4.85465e-32,-1.18662e-32) (5.51839e-34,-5.64499e-33) (-5.66765e-34,-2.6474e-34) (-4.6808e-35,4.95394e-35) 
  (-2.81088e-39,-4.03546e-40) (1.55787e-39,3.05526e-38) (3.07549e-37,-8.01782e-38) (-1.43723e-36,-2.8503e-36) (-2.393e-35,1.96523e-35) (2.29896e-34,1.76136e-34) (1.05137e-33,-2.38594e-33) (-2.22227e-32,-3.73361e-33) (1.70545e-32,1.8563e-31) (1.37747e-30,-5.18002e-31) (-6.5658e-30,-8.86812e-30) (-4.72392e-29,6.24816e-29) (4.91579e-28,1.80573e-28) (1.66191e-28,-3.27582e-27) (-1.85687e-26,4.87595e-27) (5.60919e-26,8.77014e-26) (3.32989e-25,-4.02514e-25) (-2.24382e-24,-8.91526e-25) (-7.91852e-25,1.01502e-23) (3.92377e-23,-8.09178e-24) (-6.81697e-23,-1.3092e-22) (-3.83336e-22,3.63962e-22) (1.66858e-21,7.45864e-22) (-4.27518e-22,-5.49862e-21) (-1.19434e-20,9.81131e-21) (3.75316e-20,-6.30802e-22) (-5.98437e-20,-2.36547e-20) (5.48069e-20,4.45075e-20) (-1.84502e-20,-5.93703e-20) (6.26558e-21,9.02482e-20) (-7.41218e-20,-1.0898e-19) (1.39953e-19,2.24352e-20) (-1.11574e-19,1.10639e-19) (-1.50318e-20,-1.29209e-19) (1.32675e-19,4.04009e-20) (-2.14494e-20,8.72686e-20) (-6.81991e-20,-1.90451e-20) (-8.44278e-21,-6.79192e-20) (1.11666e-21,-4.6008e-20) (-4.87194e-21,3.67577e-21) (2.02956e-21,2.23752e-20) (4.92832e-21,1.08789e-20) (1.79748e-21,1.68931e-22) (-2.11552e-22,-1.61056e-21) (-2.63446e-22,-6.47645e-22) (-4.44025e-23,-9.94093e-23) (2.23625e-23,2.34337e-23) (2.71217e-23,1.64429e-23) (1.37152e-23,-7.93732e-25) (2.75093e-24,-3.51034e-24) (-3.76795e-25,-1.20322e-24) (-2.99756e-25,-7.84555e-26) (-4.57661e-26,4.7733e-26) (4.34768e-27,1.19065e-26) (2.21703e-27,1.64608e-28) (1.63931e-28,-3.17591e-28) (-3.4614e-29,-4.00298e-29) (-6.84323e-30,2.50231e-30) (1.16877e-33,9.41104e-31) (1.08337e-31,3.80441e-32) (8.3301e-33,-1.05586e-32) (-8.24085e-34,-1.29171e-33) (-1.64986e-34,3.86827e-35) (-1.61949e-36,1.83327e-35) 
  (-7.18706e-40,3.4232e-40) (5.10287e-39,6.88712e-39) (5.9296e-38,-6.63232e-38) (-7.75182e-37,-4.41771e-37) (-2.53431e-36,8.25532e-36) (8.03258e-35,5.52802e-36) (-1.2211e-34,-7.1144e-34) (-5.6689e-33,2.52269e-33) (3.1956e-32,3.97441e-32) (2.33623e-31,-3.2398e-31) (-2.7919e-30,-1.00785e-30) (-1.23313e-30,2.08267e-29) (1.34086e-28,-3.23785e-29) (-4.38381e-28,-7.33398e-28) (-3.27311e-27,3.70145e-27) (2.4249e-26,1.06394e-26) (1.37137e-26,-1.30834e-25) (-5.89209e-25,1.21988e-25) (1.20426e-24,2.22637e-24) (7.16735e-24,-6.99826e-24) (-3.25108e-23,-1.86751e-23) (-2.93888e-23,1.34427e-22) (4.62854e-22,-1.00123e-22) (-9.58499e-22,-1.05824e-21) (-6.81483e-22,3.91164e-21) (6.58206e-21,-6.36643e-21) (-1.3659e-20,5.39258e-21) (1.52547e-20,-3.13154e-22) (-1.2061e-20,-8.21463e-21) (1.68549e-20,1.35792e-20) (-3.01822e-20,-2.91795e-21) (2.34685e-20,-2.23018e-20) (3.64647e-21,3.52446e-20) (-2.50101e-20,-1.37611e-20) (2.409e-20,-1.72982e-20) (1.4211e-20,1.48148e-20) (-1.0992e-20,1.01558e-20) (-1.23802e-20,-7.36368e-21) (-8.22184e-21,-8.10135e-21) (-1.19762e-21,2.87276e-22) (3.53599e-21,3.0177e-21) (2.67545e-21,1.08054e-21) (4.75124e-22,-2.02693e-22) (-2.61223e-22,-2.26083e-22) (-1.59153e-22,-6.39729e-23) (-3.05342e-23,-8.37907e-24) (5.88346e-24,-6.37262e-26) (6.87834e-24,-2.04041e-24) (2.09741e-24,-2.47752e-24) (-1.23176e-25,-1.0648e-24) (-2.6699e-25,-1.48228e-25) (-6.69847e-26,3.58408e-26) (-5.28072e-28,1.64145e-26) (2.78493e-27,1.53025e-27) (4.53184e-28,-3.32789e-28) (-2.00479e-29,-8.90391e-29) (-1.34492e-29,-2.29616e-30) (-9.74233e-31,1.62573e-30) (1.54212e-31,1.92747e-31) (2.87088e-32,-9.84134e-33) (1.21608e-35,-3.57256e-33) (-3.85415e-34,-1.35208e-34) (-2.826e-35,3.54163e-35) (2.69021e-36,4.10869e-36) 
  (-1.13732e-40,1.8846e-40) (2.22423e-39,8.11765e-40) (3.58096e-39,-2.42769e-38) (-2.45106e-37,1.59713e-38) (6.67306e-37,2.27505e-36) (1.9174e-35,-1.08445e-35) (-1.34575e-34,-1.43313e-34) (-9.03233e-34,1.41701e-33) (1.30737e-32,4.15953e-33) (4.06766e-33,-1.06522e-31) (-7.62507e-31,1.87482e-31) (2.76046e-30,4.71635e-30) (2.42262e-29,-2.62817e-29) (-1.97918e-28,-9.38209e-29) (-1.68649e-28,1.24049e-27) (6.53918e-27,-1.14302e-27) (-1.50708e-26,-2.89877e-26) (-1.05229e-25,1.04435e-25) (5.46558e-25,3.02554e-25) (5.68932e-25,-2.4288e-24) (-9.51258e-24,4.92317e-25) (1.35675e-23,3.28585e-23) (7.98172e-23,-9.13749e-23) (-3.60242e-22,-6.05728e-23) (5.18104e-22,8.52863e-22) (1.12224e-22,-2.17744e-21) (-1.42827e-21,2.95103e-21) (2.48761e-21,-2.12711e-21) (-3.41794e-21,3.44731e-22) (5.00309e-21,-8.08813e-22) (-4.83291e-21,4.8659e-21) (-7.85064e-22,-7.27915e-21) (6.56867e-21,4.2334e-21) (-5.58892e-21,2.71762e-21) (1.2795e-22,-6.19421e-21) (4.5883e-21,-8.40043e-22) (6.60791e-22,3.10981e-21) (-2.71176e-21,1.11985e-21) (-2.75718e-21,1.27285e-22) (-4.70624e-22,2.36901e-22) (9.14972e-22,-5.7839e-23) (6.25758e-22,-2.51353e-22) (7.85085e-23,-1.23019e-22) (-7.0681e-23,-8.49841e-25) (-3.74056e-23,1.62624e-23) (-7.328e-24,4.82448e-24) (6.30138e-25,-6.67139e-25) (6.92814e-25,-1.42914e-24) (-8.29845e-26,-7.51204e-25) (-1.99232e-25,-1.58504e-25) (-7.07417e-26,1.85566e-26) (-5.95262e-27,1.74127e-26) (2.60626e-27,3.07295e-27) (7.68431e-28,-1.71037e-28) (3.16183e-29,-1.3689e-28) (-1.83481e-29,-1.39039e-29) (-3.01046e-30,1.73401e-30) (6.9554e-32,4.81868e-31) (6.2393e-32,1.3941e-32) (4.27531e-33,-6.66669e-33) (-5.76637e-34,-7.38737e-34) (-1.01748e-34,3.46891e-35) (-7.82165e-38,1.1961e-35) (1.22787e-36,4.12357e-37) 
  (2.22412e-42,5.99996e-41) (6.27924e-40,-1.47173e-40) (-2.80541e-39,-6.05355e-39) (-5.32032e-38,4.01029e-38) (4.88662e-37,4.15009e-37) (2.70779e-36,-5.27983e-36) (-5.12668e-35,-1.22015e-35) (7.50447e-36,4.47768e-34) (3.49232e-33,-9.94726e-34) (-1.45943e-32,-2.38831e-32) (-1.38094e-31,1.50652e-31) (1.2666e-30,6.15792e-31) (1.41512e-30,-9.0058e-30) (-5.46868e-29,8.04294e-30) (1.36494e-28,2.81062e-28) (1.19286e-27,-1.12711e-27) (-6.98607e-27,-3.91958e-27) (-7.79026e-27,3.53334e-26) (1.53041e-25,-9.19515e-27) (-2.04385e-25,-5.85201e-25) (-1.95074e-24,1.42791e-24) (7.6955e-24,4.84953e-24) (2.20029e-24,-3.06585e-23) (-8.03804e-23,4.51177e-23) (2.34285e-22,7.26736e-23) (-3.25402e-22,-3.89019e-22) (2.00851e-22,6.88647e-22) (1.31795e-22,-6.88863e-22) (-5.43575e-22,5.91563e-22) (6.16703e-22,-9.85795e-22) (1.68273e-22,1.51799e-21) (-1.39795e-21,-8.51729e-22) (1.59726e-21,-5.41869e-22) (-2.15692e-22,1.32507e-21) (-1.00681e-21,-7.68231e-22) (4.26172e-22,-9.55453e-22) (6.48887e-22,2.14496e-22) (-1.29393e-22,5.64944e-22) (-4.04967e-22,4.86312e-22) (-8.30047e-23,1.62291e-22) (1.15901e-22,-1.25119e-22) (6.22616e-23,-1.39285e-22) (-3.7673e-24,-3.9377e-23) (-1.10733e-23,8.4433e-24) (-3.4656e-24,8.74449e-24) (-3.70024e-25,2.29832e-24) (3.42148e-28,-9.80828e-26) (-1.26503e-25,-3.19033e-25) (-1.38298e-25,-1.04399e-25) (-5.93437e-26,6.85789e-27) (-9.02515e-27,1.4785e-26) (1.80983e-27,4.01631e-27) (9.68785e-28,1.25287e-28) (1.13128e-28,-1.56092e-28) (-1.6215e-29,-3.06748e-29) (-5.72863e-30,3.16776e-31) (-3.02666e-31,8.19868e-31) (9.11205e-32,8.34333e-32) (1.46624e-32,-7.24581e-33) (-2.08796e-34,-2.03053e-33) (-2.35876e-34,-5.77353e-35) (-1.52114e-35,2.34442e-35) (1.91353e-36,2.46291e-36) (3.18075e-37,-1.13473e-37) 
  (9.31255e-42,1.32047e-41) (1.1974e-40,-1.25237e-40) (-1.51671e-39,-9.47979e-40) (-6.03824e-39,1.67569e-38) (1.695e-37,2.11376e-38) (-1.68641e-37,-1.56526e-36) (-1.30723e-35,4.75523e-36) (6.64105e-35,9.69293e-35) (6.15143e-34,-7.18712e-34) (-6.55777e-33,-3.05236e-33) (-8.04099e-33,5.17306e-32) (3.53971e-31,-4.83822e-32) (-9.59082e-31,-2.07875e-30) (-1.0207e-29,9.19616e-30) (6.6169e-29,3.91184e-29) (9.24355e-29,-3.89584e-28) (-1.93757e-27,1.24307e-28) (3.0043e-27,8.23254e-27) (3.04449e-26,-2.18612e-26) (-1.20875e-25,-9.52379e-26) (-2.09398e-25,5.74614e-25) (2.2974e-24,-1.46626e-25) (-4.2293e-24,-6.43234e-24) (-8.32462e-24,2.13325e-23) (5.36787e-23,-2.44387e-23) (-1.14402e-22,-1.49135e-23) (1.30383e-22,8.22719e-23) (-6.9521e-23,-1.33944e-22) (2.03999e-24,1.85344e-22) (-7.83397e-23,-2.49822e-22) (2.8384e-22,1.78656e-22) (-3.37354e-22,1.29284e-22) (1.18251e-22,-3.36419e-22) (2.05197e-22,2.01452e-22) (-2.42377e-22,7.59273e-23) (-1.17837e-22,-1.97948e-22) (1.11945e-22,-9.81319e-23) (7.74177e-23,8.05589e-23) (1.97604e-23,1.38181e-22) (1.37607e-23,5.20331e-23) (1.82777e-25,-2.93667e-23) (-1.14431e-23,-3.13963e-23) (-7.32764e-24,-7.16592e-24) (-8.20761e-25,2.53246e-24) (8.14327e-25,1.94034e-24) (3.61817e-25,4.71243e-25) (5.77075e-27,1.24546e-27) (-6.73956e-26,-2.58221e-26) (-3.85388e-26,6.57206e-27) (-8.54625e-27,1.08905e-26) (8.89671e-28,3.95897e-27) (9.63409e-28,3.98367e-28) (1.91414e-28,-1.34705e-28) (-4.68965e-30,-4.64344e-29) (-7.90295e-30,-3.05069e-30) (-1.02268e-30,9.75373e-31) (7.32222e-32,2.04547e-31) (3.09377e-32,1.62696e-33) (1.72486e-33,-3.75699e-33) (-3.64646e-34,-3.70412e-34) (-5.65246e-35,2.59108e-35) (6.59808e-37,7.1492e-36) (7.79974e-37,1.93289e-37) (4.63624e-38,-7.3688e-38) 
  (3.98219e-42,1.599e-42) (8.5617e-42,-4.51185e-41) (-4.72808e-40,8.39928e-42) (1.078e-39,4.56939e-39) (4.02963e-38,-1.9705e-38) (-2.61259e-37,-3.18014e-37) (-2.15977e-36,2.90134e-36) (2.81218e-35,1.14443e-35) (2.97092e-35,-2.40859e-34) (-1.81974e-33,2.76458e-34) (5.54208e-33,1.19847e-32) (6.68912e-32,-5.90736e-32) (-4.8229e-31,-2.96796e-31) (-8.39692e-31,3.25844e-30) (1.86326e-29,-8.89798e-31) (-3.25223e-29,-9.08532e-29) (-3.75399e-28,2.76062e-28) (1.66924e-27,1.29208e-27) (3.4473e-27,-8.46641e-27) (-3.80004e-26,-3.64638e-27) (3.81156e-26,1.49035e-25) (4.41146e-25,-3.70108e-25) (-1.80297e-24,-6.14787e-25) (1.77717e-24,5.3032e-24) (5.57176e-24,-1.27083e-23) (-2.10516e-23,1.47284e-23) (3.22711e-23,-4.88138e-24) (-2.98054e-23,-1.34017e-23) (2.9828e-23,2.95967e-23) (-5.35044e-23,-2.22457e-23) (6.85006e-23,-2.43773e-23) (-2.28201e-23,7.51857e-23) (-4.02594e-23,-6.2035e-23) (6.0022e-23,-1.07638e-23) (-1.44927e-23,4.80603e-23) (-4.94531e-23,-4.29902e-24) (-5.69214e-24,-3.2209e-23) (2.07462e-23,-4.94094e-24) (2.4728e-23,1.63923e-23) (1.2321e-23,7.45594e-24) (-2.8598e-24,-3.48595e-24) (-6.37253e-24,-3.08843e-24) (-2.54222e-24,-1.27704e-25) (1.06499e-25,4.96213e-25) (4.19178e-25,1.81138e-25) (1.45443e-25,1.63938e-26) (7.48803e-27,-1.70867e-27) (-1.31748e-26,6.5468e-27) (-4.78976e-27,7.23101e-27) (4.04595e-28,3.14103e-27) (7.87516e-28,5.13404e-28) (2.27826e-28,-8.72551e-29) (1.17097e-29,-5.41904e-29) (-8.25627e-30,-7.52717e-30) (-1.92089e-30,7.02442e-31) (-3.43097e-32,3.4244e-31) (4.61466e-32,2.68437e-32) (6.16328e-33,-4.57983e-33) (-2.59126e-34,-9.99734e-34) (-1.2993e-34,-1.51087e-35) (-7.11493e-36,1.40375e-35) (1.25713e-36,1.32068e-36) (1.86448e-37,-8.43606e-38) (-2.32683e-39,-2.20735e-38) 
  (1.10445e-42,-2.13291e-43) (-4.52255e-42,-1.11269e-41) (-1.02306e-40,6.88867e-41) (8.82238e-40,8.43245e-40) (5.95145e-39,-9.97292e-39) (-1.01209e-37,-3.16771e-38) (-5.40843e-38,9.25175e-37) (7.57993e-36,-1.51109e-36) (-2.73384e-35,-5.48928e-35) (-3.417e-34,3.09934e-34) (2.7945e-33,1.71745e-33) (5.66842e-33,-2.12157e-32) (-1.37962e-31,4.60057e-33) (2.63442e-31,7.68704e-31) (3.62323e-30,-2.61659e-30) (-1.82388e-29,-1.40146e-29) (-4.03647e-29,1.03357e-28) (5.04085e-28,5.07059e-29) (-3.88553e-28,-2.19267e-27) (-8.37367e-27,4.38951e-27) (2.91064e-26,2.50228e-26) (3.25582e-26,-1.38528e-25) (-4.38812e-25,1.54889e-25) (1.14734e-24,6.95783e-25) (-9.99735e-25,-3.03544e-24) (-1.25458e-24,5.46583e-24) (4.49628e-24,-5.14014e-24) (-6.87783e-24,1.80717e-24) (9.34162e-24,-1.68634e-25) (-1.11543e-23,5.91472e-24) (4.92051e-24,-1.47762e-23) (9.67468e-24,1.37537e-23) (-1.50344e-23,-1.08301e-24) (5.47314e-24,-1.15466e-23) (6.35756e-24,7.50925e-24) (-6.8542e-24,7.88824e-24) (-6.65401e-24,-2.7221e-24) (1.00471e-24,-4.01739e-24) (5.86442e-24,-1.60136e-24) (3.49091e-24,-8.60807e-25) (-5.38491e-25,-1.93099e-25) (-1.37743e-24,4.52475e-25) (-4.69719e-25,3.86225e-25) (6.21382e-26,8.12395e-26) (9.03477e-26,-3.26976e-26) (2.70663e-26,-2.20301e-26) (1.74329e-27,-2.65236e-27) (-8.01375e-28,2.77749e-27) (4.3708e-28,1.83937e-27) (5.70787e-28,4.30551e-28) (2.11213e-28,-4.22071e-29) (2.42914e-29,-5.09725e-29) (-6.61686e-30,-1.1172e-29) (-2.64506e-30,-1.39973e-32) (-2.3348e-31,4.29013e-31) (4.76176e-32,6.78353e-32) (1.27703e-32,-2.27151e-33) (4.4256e-34,-1.82882e-33) (-2.06018e-34,-1.50397e-34) (-2.74997e-35,1.73989e-35) (8.01007e-37,3.85583e-36) (4.53427e-37,6.39031e-38) (2.368e-38,-4.57708e-38) (-3.9044e-39,-4.01101e-39) 
  (2.10688e-43,-2.00864e-43) (-2.53645e-42,-1.78307e-42) (-1.24962e-41,2.91785e-41) (3.07463e-40,5.83417e-41) (-1.16e-40,-2.9631e-39) (-2.59231e-38,7.33637e-39) (1.16831e-37,2.02811e-37) (1.37902e-36,-1.36304e-36) (-1.32156e-35,-7.64605e-36) (-2.80705e-35,1.10403e-34) (8.02306e-34,-2.75298e-35) (-1.69231e-33,-5.04912e-33) (-2.708e-32,1.91598e-32) (1.52738e-31,1.19011e-31) (3.84929e-31,-9.85792e-31) (-5.40942e-30,-4.81465e-31) (4.87696e-30,2.58153e-29) (1.08955e-28,-5.34584e-29) (-3.65699e-28,-4.00088e-28) (-1.12018e-27,2.04715e-27) (9.44545e-27,8.50823e-28) (-1.41042e-26,-3.17399e-26) (-5.92046e-26,9.52238e-26) (3.11844e-25,-5.12107e-26) (-6.25144e-25,-3.59167e-25) (5.7892e-25,1.05275e-24) (3.77094e-26,-1.41707e-24) (-8.96893e-25,1.26166e-24) (1.36495e-24,-1.51216e-24) (-5.23564e-25,2.66124e-24) (-1.83035e-24,-2.74246e-24) (3.53277e-24,1.82053e-25) (-1.96999e-24,2.29816e-24) (-1.27873e-24,-2.31048e-24) (1.90727e-24,-2.83627e-25) (4.81439e-25,2.09363e-24) (-1.29364e-24,8.85363e-25) (-6.52271e-25,-5.37231e-25) (5.12147e-25,-1.08556e-24) (4.3184e-25,-7.32757e-25) (-6.11792e-26,-2.9551e-26) (-1.34106e-25,2.52677e-25) (-1.88937e-26,1.38893e-25) (2.01903e-26,1.10125e-26) (9.06562e-27,-1.73644e-26) (7.98932e-28,-8.02996e-27) (-2.03948e-28,-1.00038e-27) (2.85255e-28,4.62114e-28) (3.51594e-28,2.00041e-28) (1.57352e-28,-2.42779e-29) (2.73752e-29,-4.03933e-29) (-4.04288e-30,-1.2279e-29) (-2.88534e-30,-8.48118e-31) (-4.60907e-31,4.13817e-31) (2.58852e-32,1.12453e-31) (1.91572e-32,4.77356e-33) (1.98196e-33,-2.40526e-33) (-2.02243e-34,-4.08665e-34) (-6.21906e-35,3.64645e-36) (-2.55169e-36,7.58764e-36) (7.51714e-37,6.20286e-37) (9.80586e-38,-5.76537e-38) (-2.44721e-39,-1.26008e-38) (-1.38462e-39,-1.8314e-40) 
  (1.76881e-44,-7.22488e-44) (-7.89404e-43,-3.32188e-44) (1.34661e-42,7.94908e-42) (7.33282e-41,-2.98741e-41) (-4.31262e-40,-6.09761e-40) (-4.43248e-39,5.08975e-39) (5.20186e-38,2.62741e-38) (9.95095e-38,-4.6901e-37) (-3.73993e-36,2.20415e-37) (9.1135e-36,2.61802e-35) (1.57826e-34,-1.12187e-34) (-1.00156e-33,-7.8591e-34) (-2.88726e-33,7.31458e-33) (4.53934e-32,3.99086e-33) (-4.8158e-32,-2.43262e-31) (-1.13352e-30,5.78382e-31) (4.18568e-30,4.57201e-30) (1.53882e-29,-2.46413e-29) (-1.27368e-28,-3.38339e-29) (5.52053e-29,5.70171e-28) (1.98805e-27,-1.19055e-27) (-7.35844e-27,-3.99007e-27) (3.34277e-27,2.64162e-26) (4.68235e-26,-5.60643e-26) (-1.55985e-25,3.29799e-26) (2.37988e-25,8.59754e-26) (-1.7918e-25,-2.31779e-25) (3.2697e-26,3.33557e-25) (-4.40682e-26,-4.33616e-25) (3.70852e-25,4.39657e-25) (-6.88199e-25,-4.88705e-26) (4.79823e-25,-5.51454e-25) (1.40927e-25,5.83924e-25) (-5.33528e-25,-6.35946e-26) (1.45416e-25,-3.5211e-25) (3.974e-25,1.68007e-25) (4.63455e-28,3.36863e-25) (-1.66663e-25,7.66896e-26) (-9.69005e-26,-2.06476e-25) (-5.15225e-26,-1.8529e-25) (-1.87738e-26,-1.44884e-26) (1.45266e-26,5.21821e-26) (1.80994e-26,2.5465e-26) (5.64351e-27,1.14271e-28) (-9.36446e-28,-3.75086e-27) (-1.14377e-27,-1.40556e-27) (-2.42572e-28,-1.60517e-28) (9.48363e-29,1.64339e-29) (8.0947e-29,-2.553e-29) (2.01828e-29,-2.85445e-29) (-2.01422e-30,-1.07413e-29) (-2.58706e-30,-1.37137e-30) (-6.15262e-31,3.10114e-31) (-1.42392e-32,1.42788e-31) (2.20002e-32,1.56098e-32) (4.14232e-33,-2.11967e-33) (-1.40373e-35,-7.40672e-34) (-1.00166e-34,-4.37312e-35) (-1.10089e-35,1.02612e-35) (6.866e-37,1.82274e-36) (2.38562e-37,2.77797e-39) (1.00092e-38,-2.61057e-38) (-2.40171e-39,-2.0591e-39) (-2.96431e-40,1.7627e-40) 
  (-6.04119e-45,-1.77723e-44) (-1.71784e-43,1.00062e-43) (1.36197e-42,1.49373e-42) (1.1331e-41,-1.62009e-41) (-1.72379e-40,-6.87375e-41) (-2.30411e-40,1.65168e-39) (1.42188e-38,-1.60002e-39) (-4.25085e-38,-1.08876e-37) (-7.26273e-37,5.41963e-37) (5.27975e-36,4.04257e-36) (1.6715e-35,-4.29068e-35) (-2.99082e-34,-2.59084e-35) (3.63697e-34,1.80394e-33) (9.39911e-33,-4.90811e-33) (-3.95637e-32,-4.18583e-32) (-1.53503e-31,2.53751e-31) (1.40427e-30,4.00354e-31) (-4.48039e-33,-6.95262e-30) (-3.03576e-29,1.00119e-29) (9.03268e-29,1.06388e-28) (2.14535e-28,-5.1672e-28) (-1.96417e-27,3.27874e-28) (4.52847e-27,4.27389e-27) (-3.2254e-28,-1.65667e-26) (-2.05127e-26,2.7847e-26) (4.89978e-26,-1.88419e-26) (-5.88288e-26,-1.38629e-26) (5.31921e-26,4.8228e-26) (-7.46791e-26,-5.3123e-26) (1.20467e-25,-3.54775e-27) (-9.50931e-26,1.06317e-25) (-2.82596e-26,-1.45611e-25) (1.09873e-25,4.35574e-26) (-7.26779e-26,7.92148e-26) (-4.59411e-26,-6.08843e-26) (7.21695e-26,-4.44753e-26) (5.823e-26,4.0687e-26) (-2.57957e-27,4.14145e-26) (-4.05649e-26,-9.42413e-27) (-3.68654e-26,-1.96663e-26) (-8.44334e-27,-1.26692e-27) (8.33282e-27,5.11657e-27) (6.6129e-27,1.31678e-27) (1.21222e-27,-7.33481e-28) (-5.99498e-28,-4.30753e-28) (-3.93125e-28,-4.39821e-29) (-7.52235e-29,1.523e-29) (1.19905e-29,-1.01664e-29) (7.41268e-30,-1.57928e-29) (-1.42784e-30,-7.42968e-30) (-1.99479e-30,-1.36863e-30) (-6.30512e-31,1.81604e-31) (-5.33508e-32,1.46765e-31) (1.97257e-32,2.63181e-32) (6.20073e-33,-7.04679e-34) (4.00582e-34,-1.00866e-33) (-1.16144e-34,-1.29867e-34) (-2.48333e-35,7.42511e-36) (-4.53157e-37,3.56816e-36) (4.06061e-37,2.34386e-37) (4.53355e-38,-3.58301e-38) (-2.0668e-39,-6.47912e-39) (-7.71128e-40,-2.8846e-41) (-3.0137e-41,7.87262e-41) 
  (-3.64824e-45,-2.92969e-45) (-2.25867e-44,4.3931e-44) (4.83438e-43,1.2907e-43) (1.82586e-43,-4.86874e-42) (-4.4632e-41,8.84455e-42) (1.72595e-40,3.68025e-40) (2.67007e-39,-2.20795e-39) (-2.28922e-38,-1.62884e-38) (-7.39166e-38,2.03086e-37) (1.56856e-36,1.15119e-37) (-2.21881e-36,-1.05698e-35) (-6.16895e-35,3.27921e-35) (2.95839e-34,3.05843e-34) (1.22798e-33,-2.11204e-33) (-1.28456e-32,-3.38941e-33) (4.17907e-34,6.88944e-32) (3.31155e-31,-9.28543e-32) (-8.89548e-31,-1.40511e-30) (-4.76508e-30,6.07717e-30) (3.26433e-29,8.31972e-30) (-3.32219e-29,-1.29209e-28) (-3.14124e-28,3.46187e-28) (1.43038e-27,8.94873e-29) (-2.47876e-27,-2.73273e-27) (6.58209e-28,7.33783e-27) (5.13159e-27,-9.44748e-27) (-1.12137e-26,5.43453e-27) (1.51565e-26,-3.11855e-28) (-1.83981e-26,4.64418e-27) (1.48822e-26,-2.00437e-26) (5.27941e-27,2.86368e-26) (-2.63786e-26,-1.3338e-26) (1.92381e-26,-1.28427e-26) (4.35249e-27,2.06854e-26) (-1.53783e-26,1.69098e-27) (8.94826e-28,-1.63114e-26) (1.38179e-26,-4.91433e-27) (7.76733e-27,5.40781e-27) (-5.52593e-27,4.77834e-27) (-8.29122e-27,2.79121e-27) (-2.15698e-27,1.29449e-27) (1.63862e-27,-2.94595e-28) (1.19404e-27,-7.50346e-28) (1.34516e-28,-3.21955e-28) (-1.36367e-28,6.50397e-30) (-6.64093e-29,5.14217e-29) (-1.06308e-29,1.59278e-29) (-1.9039e-31,-2.25506e-30) (-1.34299e-30,-3.24143e-30) (-1.35611e-30,-8.73644e-31) (-5.20051e-31,9.78374e-32) (-7.22628e-32,1.26255e-31) (1.39297e-32,3.21308e-32) (7.33592e-33,1.35241e-33) (9.47198e-34,-1.06995e-33) (-8.45797e-35,-2.35845e-34) (-4.02209e-35,-5.17182e-36) (-3.31078e-36,5.10282e-36) (4.59314e-37,7.15996e-37) (1.10144e-37,-1.8445e-38) (3.01295e-39,-1.35188e-38) (-1.36497e-39,-9.04519e-40) (-1.49993e-40,1.1057e-40) (6.10687e-42,1.94647e-41) 
  (-1.14506e-45,-1.27816e-46) (1.1211e-45,1.20704e-44) (1.16508e-43,-3.71766e-44) (-6.0385e-43,-1.01985e-42) (-7.90404e-42,7.66284e-42) (8.30235e-41,5.15963e-41) (2.46208e-40,-7.90045e-40) (-6.65523e-39,-2.64973e-40) (1.15654e-38,4.9497e-38) (3.21254e-37,-1.77236e-37) (-1.76071e-36,-1.77425e-36) (-7.86796e-36,1.39988e-35) (9.45902e-35,2.29612e-35) (-1.65871e-35,-5.58095e-34) (-2.92113e-33,8.76951e-34) (8.39581e-33,1.36052e-32) (5.49095e-32,-5.96058e-32) (-3.60066e-31,-1.67613e-31) (-1.25801e-31,1.85039e-30) (7.48016e-30,-2.9616e-30) (-2.46753e-29,-1.94328e-29) (-6.75377e-30,1.08029e-28) (2.61024e-28,-1.92829e-28) (-8.01193e-28,-9.33311e-29) (1.11704e-27,1.06383e-27) (-4.35635e-28,-2.13489e-27) (-1.07054e-27,2.33142e-27) (2.19864e-27,-2.2509e-27) (-1.66902e-27,3.49957e-27) (-1.34336e-27,-4.93307e-27) (5.2126e-27,2.69038e-27) (-5.21757e-27,2.50613e-27) (4.21433e-29,-4.51334e-27) (3.74993e-27,1.62152e-27) (-1.34667e-27,2.86044e-27) (-2.47333e-27,-1.86815e-27) (8.21602e-28,-2.8455e-27) (1.98205e-27,-7.7425e-28) (1.76451e-28,1.22673e-27) (-7.30338e-28,1.61006e-27) (-1.85039e-28,6.30887e-28) (1.70249e-28,-2.0008e-28) (7.14685e-29,-2.76781e-28) (-2.28474e-29,-7.98801e-29) (-1.92571e-29,1.53102e-29) (-2.56023e-30,1.71589e-29) (8.70498e-31,4.48604e-30) (-2.63009e-31,-7.11285e-32) (-6.50356e-31,-2.29248e-31) (-3.29064e-31,8.05347e-32) (-6.40236e-32,9.47552e-32) (8.00067e-33,3.089e-32) (7.15366e-33,3.03729e-33) (1.41353e-33,-8.9737e-34) (-3.6054e-36,-3.23876e-34) (-5.02121e-35,-2.75286e-35) (-7.7747e-36,5.18139e-36) (1.85503e-37,1.40066e-36) (1.90155e-37,5.90823e-38) (1.7223e-38,-1.99132e-38) (-1.47542e-39,-2.93614e-39) (-3.88631e-40,3.64418e-41) (-1.152e-41,4.30426e-41) (4.0457e-42,2.74504e-42) 
  (-2.52003e-46,1.2274e-46) (1.79976e-45,2.3227e-45) (1.88557e-44,-2.27077e-44) (-2.54407e-43,-1.27629e-43) (-5.93046e-43,2.56098e-42) (2.31891e-41,-4.41166e-43) (-5.27893e-41,-1.87691e-40) (-1.33836e-39,7.96552e-40) (8.50457e-39,8.16938e-39) (3.9953e-38,-7.44051e-38) (-5.57556e-37,-1.24201e-37) (1.91015e-37,3.64427e-36) (2.09492e-35,-6.9199e-36) (-6.94388e-35,-1.0614e-34) (-4.68186e-34,5.18352e-34) (3.30544e-33,1.68775e-33) (3.54968e-33,-1.87686e-32) (-9.35867e-32,1.35358e-32) (2.26921e-31,3.79282e-31) (1.00696e-30,-1.61027e-30) (-7.29877e-30,-6.40365e-32) (1.43087e-29,2.01474e-29) (1.66153e-29,-7.03423e-29) (-1.42769e-28,9.8108e-29) (3.17549e-28,1.44146e-29) (-3.41519e-28,-2.74279e-28) (1.3985e-28,5.07216e-28) (-1.37722e-29,-6.41055e-28) (3.37127e-28,7.07382e-28) (-9.53459e-28,-4.02622e-28) (1.05634e-27,-4.91885e-28) (-2.2189e-28,1.0926e-27) (-7.23536e-28,-4.9922e-28) (6.60169e-28,-4.09889e-28) (3.45545e-28,5.45457e-28) (-5.47186e-28,1.99289e-28) (-3.62297e-28,-4.59611e-28) (1.15273e-28,-4.51967e-28) (1.9717e-28,6.95186e-29) (1.34529e-28,3.17643e-28) (7.38027e-29,1.40547e-28) (4.19641e-30,-3.72532e-29) (-2.70027e-29,-4.9207e-29) (-1.58452e-29,-1.06232e-29) (-1.46201e-30,4.14915e-30) (1.99192e-30,2.86056e-30) (8.65812e-31,5.94239e-31) (1.9741e-33,4.77945e-32) (-1.15386e-31,6.4696e-32) (-3.44543e-32,6.09946e-32) (4.84773e-33,2.39241e-32) (5.93499e-33,3.56717e-33) (1.59678e-33,-6.0321e-34) (9.36801e-35,-3.59969e-34) (-4.95202e-35,-5.32001e-35) (-1.26286e-35,2.90429e-36) (-5.57682e-37,2.05695e-36) (2.4222e-37,2.16528e-37) (4.24929e-38,-1.79834e-38) (1.16343e-40,-6.14333e-39) (-7.0536e-40,-3.1327e-40) (-6.58742e-41,6.44197e-41) (4.24565e-42,9.66056e-42) (1.15728e-42,-8.76664e-44) 
  (-3.54555e-47,5.72962e-47) (6.61892e-46,2.38524e-46) (8.76697e-46,-6.97983e-45) (-6.7107e-44,7.09039e-45) (2.09303e-43,5.83114e-43) (4.5042e-42,-3.03309e-42) (-3.40061e-41,-2.99618e-41) (-1.59452e-40,3.2198e-40) (2.64959e-39,5.16991e-40) (-1.47019e-39,-1.91344e-38) (-1.21388e-37,4.36633e-38) (4.70395e-37,6.72897e-37) (3.20523e-36,-3.79132e-36) (-2.58717e-35,-1.24401e-35) (-3.07414e-35,1.56934e-34) (8.60142e-34,-6.49398e-35) (-1.65738e-33,-4.18221e-33) (-1.6658e-32,1.4982e-32) (9.54974e-32,4.20719e-32) (-3.7038e-32,-4.41347e-31) (-1.32722e-30,1.02025e-30) (5.36184e-30,1.47371e-30) (-7.22081e-30,-1.40896e-29) (-9.10596e-30,3.5414e-29) (5.07991e-29,-3.98426e-29) (-8.75196e-29,1.07203e-30) (8.90861e-29,5.95218e-29) (-9.50379e-29,-8.61285e-29) (1.52937e-28,3.53609e-29) (-1.8106e-28,1.00305e-28) (5.02077e-29,-2.22539e-28) (1.41184e-28,1.57566e-28) (-1.59091e-28,6.21008e-29) (5.82789e-30,-1.45686e-28) (1.30774e-28,2.31918e-30) (-2.24974e-29,1.0677e-28) (-1.13157e-28,5.66075e-30) (-6.22368e-29,-7.73508e-29) (2.48683e-29,-2.80592e-29) (6.1305e-29,2.13977e-29) (3.4466e-29,1.08777e-29) (-1.12264e-30,-4.82148e-30) (-1.01237e-29,-3.34566e-30) (-4.19394e-30,5.39795e-31) (1.22097e-31,8.02055e-31) (6.65258e-31,1.45328e-31) (2.29911e-31,-4.02616e-32) (1.76074e-32,1.93108e-33) (-4.77527e-33,2.42845e-32) (4.31507e-33,1.35922e-32) (4.32388e-33,2.78985e-33) (1.4446e-33,-3.50524e-34) (1.59501e-34,-3.35027e-34) (-3.91093e-35,-7.18405e-35) (-1.6096e-35,-1.29166e-36) (-1.67453e-36,2.3724e-36) (2.11938e-37,4.32234e-37) (7.39611e-38,1.28409e-39) (4.76077e-39,-9.45573e-39) (-8.9007e-40,-1.1062e-39) (-1.72921e-40,4.8133e-41) (-2.44492e-42,2.14002e-41) (2.19642e-42,1.14202e-42) (1.99974e-43,-1.85782e-43) 
  (1.32785e-49,1.60032e-47) (1.6244e-46,-3.61278e-47) (-7.08335e-46,-1.49659e-45) (-1.23379e-44,9.86216e-45) (1.14253e-43,8.7843e-44) (4.95952e-43,-1.15245e-42) (-1.02783e-41,-1.55696e-42) (9.06702e-42,8.12892e-41) (5.67476e-40,-2.23828e-40) (-2.57543e-39,-3.45354e-39) (-1.78453e-38,2.26352e-38) (1.67973e-37,7.30955e-38) (1.76237e-37,-1.09764e-36) (-6.46291e-36,5.82011e-37) (1.24558e-35,3.44767e-35) (1.62484e-34,-1.17766e-34) (-8.59799e-34,-6.149e-34) (-1.25137e-33,5.12237e-33) (2.38418e-32,-5.09854e-33) (-6.82531e-32,-7.57897e-32) (-9.22154e-32,3.67466e-31) (1.12514e-30,-5.04221e-31) (-3.15541e-30,-1.29548e-30) (3.39454e-30,6.79051e-30) (2.57912e-30,-1.2684e-29) (-1.33158e-29,1.12128e-29) (2.13827e-29,-2.97998e-30) (-2.50875e-29,2.37611e-30) (2.43067e-29,-1.95812e-29) (-6.49869e-30,4.03476e-29) (-2.81102e-29,-3.38564e-29) (3.9436e-29,-3.9726e-30) (-7.37389e-30,3.22021e-29) (-2.20206e-29,-1.57835e-29) (1.50456e-29,-2.13632e-29) (1.50268e-29,1.40042e-29) (-1.14307e-29,1.82581e-29) (-2.0497e-29,4.21398e-31) (-3.56406e-30,-6.75375e-30) (1.02744e-29,-5.73792e-30) (6.946e-30,-3.64953e-30) (-1.82336e-31,-8.79503e-31) (-1.7834e-30,8.01497e-31) (-5.93488e-31,6.85279e-31) (9.13274e-32,1.33268e-31) (1.12082e-31,-6.43425e-32) (2.94702e-32,-4.07959e-32) (3.61699e-33,-4.42594e-33) (2.89088e-33,3.47137e-33) (2.59062e-33,1.2064e-33) (1.04322e-33,-2.43021e-34) (1.65079e-34,-2.6907e-34) (-2.53874e-35,-7.56991e-35) (-1.69223e-35,-5.54388e-36) (-2.7983e-36,2.18843e-36) (7.59078e-38,6.3999e-37) (9.95319e-38,4.11269e-38) (1.27878e-38,-1.07083e-38) (-5.71694e-40,-2.33645e-39) (-3.18782e-40,-6.27746e-41) (-2.36028e-41,3.39419e-41) (2.69637e-42,4.196e-42) (5.6399e-43,-1.14047e-43) (9.36669e-45,-6.29178e-44) 
  (2.02586e-48,3.16282e-48) (2.75732e-47,-2.7413e-47) (-3.25479e-46,-2.05398e-46) (-1.17883e-45,3.45457e-45) (3.29676e-44,2.86112e-45) (-4.64236e-44,-2.82292e-43) (-2.1501e-42,9.5625e-43) (1.15277e-41,1.43156e-41) (8.04219e-41,-1.09861e-40) (-8.90813e-40,-3.47979e-40) (-7.46783e-40,6.33785e-39) (4.02731e-38,-5.34164e-39) (-9.13555e-38,-2.30936e-37) (-1.19096e-36,8.58377e-37) (6.53512e-36,5.30831e-36) (1.75341e-35,-4.32631e-35) (-2.4717e-34,-9.57165e-36) (4.43764e-34,1.14804e-33) (3.73992e-33,-4.21063e-33) (-2.28051e-32,-4.19938e-33) (3.51627e-32,7.69377e-32) (1.18611e-31,-2.41791e-31) (-6.86417e-31,2.26932e-31) (1.43235e-30,5.96369e-31) (-1.22864e-30,-2.25285e-30) (-6.22159e-31,3.3908e-30) (2.73025e-30,-3.31138e-30) (-2.86194e-30,3.94113e-30) (-1.01484e-31,-6.16437e-30) (5.39831e-30,5.84987e-30) (-8.35585e-30,3.32522e-31) (3.64922e-30,-6.38041e-30) (4.30056e-30,4.66654e-30) (-4.65168e-30,1.86616e-30) (-1.76838e-30,-4.81573e-30) (3.7477e-30,-1.10044e-30) (1.62127e-30,3.69694e-30) (-2.46644e-30,3.28599e-30) (-1.71437e-30,9.06461e-32) (4.07686e-31,-2.00574e-30) (4.70475e-31,-1.56585e-30) (-1.08873e-31,-2.35883e-31) (-1.40752e-31,3.15032e-31) (4.01199e-33,1.88264e-31) (3.07416e-32,1.66833e-32) (7.67577e-33,-2.25364e-32) (-1.50257e-33,-1.04396e-32) (-3.04103e-34,-1.56254e-33) (8.06459e-34,-3.66618e-35) (5.1954e-34,-2.19028e-34) (1.12378e-34,-1.89322e-34) (-1.54761e-35,-6.44767e-35) (-1.51121e-35,-7.80101e-36) (-3.46995e-36,1.64063e-36) (-1.23823e-37,7.63951e-37) (1.06748e-37,9.31502e-38) (2.25485e-38,-7.816e-39) (5.81753e-40,-3.67934e-39) (-4.39908e-40,-3.15433e-40) (-6.43877e-41,3.57367e-41) (8.13061e-43,9.39647e-42) (1.08872e-42,3.5186e-43) (8.44022e-44,-1.02176e-43) (-7.40297e-45,-1.26908e-44) 
  (7.87739e-49,3.71707e-49) (2.01047e-48,-8.74592e-48) (-8.83468e-47,1.19274e-49) (1.95472e-46,8.09555e-46) (6.6528e-45,-3.46333e-45) (-4.2907e-44,-4.80073e-44) (-2.91417e-43,4.37677e-43) (3.85744e-42,1.32569e-42) (2.25086e-42,-2.99544e-41) (-2.06924e-40,3.71558e-41) (5.78106e-40,1.2783e-39) (7.0578e-39,-5.54957e-39) (-4.37188e-38,-3.41748e-38) (-1.33383e-37,3.05013e-37) (1.91912e-36,2.61844e-37) (-1.96264e-36,-1.06615e-35) (-4.89541e-35,3.02376e-35) (2.37357e-34,1.56953e-34) (1.09117e-34,-1.28073e-33) (-4.61836e-33,2.39887e-33) (1.66703e-32,8.32094e-33) (-1.38084e-32,-5.62766e-32) (-7.78118e-32,1.29162e-31) (2.97067e-31,-9.68118e-32) (-4.68688e-31,-1.85137e-31) (3.33338e-31,5.9193e-31) (-5.76516e-32,-8.377e-31) (2.18651e-31,9.02168e-31) (-9.67114e-31,-7.26238e-31) (1.5236e-30,-1.21558e-31) (-8.96292e-31,1.28418e-30) (-5.78183e-31,-1.22352e-30) (1.19558e-30,-1.68321e-31) (-1.59847e-31,9.14744e-31) (-9.55322e-31,-2.52602e-31) (1.86381e-31,-7.27631e-31) (7.38272e-31,1.28174e-31) (2.05491e-31,7.72896e-31) (-1.80606e-31,3.50301e-31) (-2.15213e-31,-2.63253e-31) (-1.59635e-31,-2.86823e-31) (-6.09534e-32,-4.08394e-32) (1.64705e-32,5.59808e-32) (2.61173e-32,2.75303e-32) (7.89581e-33,-3.1058e-34) (-1.54933e-33,-3.96147e-33) (-1.69548e-33,-1.32408e-33) (-3.4525e-34,-2.09409e-34) (7.55409e-35,-1.21149e-34) (3.53313e-35,-1.03718e-34) (-1.21477e-35,-4.30002e-35) (-1.17756e-35,-7.15054e-36) (-3.42905e-36,1.04963e-36) (-2.94924e-37,7.64273e-37) (9.26717e-38,1.38906e-37) (3.08458e-38,-6.27997e-40) (2.55389e-39,-4.57448e-39) (-4.39446e-40,-6.97215e-40) (-1.20197e-40,1.07277e-41) (-5.83517e-42,1.54704e-41) (1.50288e-42,1.51164e-42) (2.41833e-43,-9.56425e-44) (2.31653e-46,-3.02498e-44) (-3.14176e-45,-1.20155e-45) 
  (1.98199e-49,-2.34934e-50) (-6.72391e-49,-1.93233e-48) (-1.69277e-47,1.07022e-47) (1.34626e-46,1.30657e-46) (8.44381e-46,-1.45027e-45) (-1.37532e-44,-3.93838e-45) (-3.18033e-45,1.15985e-43) (8.72091e-43,-1.99279e-43) (-2.99625e-42,-5.83482e-42) (-3.44933e-41,3.02038e-41) (2.51168e-40,1.76564e-40) (7.29816e-40,-1.84369e-39) (-1.23131e-38,-1.68246e-39) (9.37724e-39,7.51208e-38) (4.07394e-37,-1.81e-37) (-1.72586e-36,-1.82033e-36) (-5.36381e-36,1.21529e-35) (6.50356e-35,-2.73508e-36) (-1.54639e-34,-2.45056e-34) (-4.75851e-34,1.0501e-33) (3.94954e-33,-8.84592e-34) (-9.91622e-33,-7.24429e-33) (5.13948e-33,3.05337e-32) (3.24283e-32,-5.29181e-32) (-9.33264e-32,3.0483e-32) (1.24655e-31,4.63677e-32) (-1.20436e-31,-1.07454e-31) (1.57582e-31,7.61247e-32) (-2.2718e-31,6.16696e-32) (1.59709e-31,-2.41047e-31) (9.03178e-32,2.74722e-31) (-2.44912e-31,-3.93921e-32) (1.02253e-31,-2.02694e-31) (1.30281e-31,1.14106e-31) (-1.42655e-31,1.20383e-31) (-1.01813e-31,-1.04054e-31) (9.3881e-32,-1.01914e-31) (1.39061e-31,5.97054e-32) (4.20019e-32,7.77526e-32) (-5.36388e-32,2.28779e-33) (-6.15034e-32,-1.62913e-32) (-1.85864e-32,1.54114e-33) (7.68763e-33,5.43982e-33) (7.4052e-33,5.48878e-34) (1.43326e-33,-1.06453e-33) (-6.37795e-34,-3.70014e-34) (-4.25317e-34,4.16391e-35) (-9.26171e-35,2.52953e-35) (-1.1488e-35,-2.28613e-35) (-1.05347e-35,-1.8159e-35) (-7.9473e-36,-4.12932e-36) (-2.7448e-36,6.94005e-37) (-3.57017e-37,6.57999e-37) (6.66645e-38,1.59797e-37) (3.47385e-38,8.16372e-39) (4.82101e-39,-4.58919e-39) (-2.50022e-40,-1.11183e-39) (-1.73278e-40,-5.11152e-41) (-1.85234e-41,1.91648e-41) (1.24399e-42,3.46138e-42) (4.75401e-43,4.28514e-44) (2.82263e-44,-5.13238e-44) (-4.28794e-45,-5.33423e-45) (-7.26166e-46,2.35682e-46) 
  (3.52696e-50,-2.82438e-50) (-3.59116e-49,-2.88646e-49) (-1.93763e-48,4.04278e-48) (4.08091e-47,8.69638e-48) (-1.20705e-47,-3.70526e-46) (-3.01766e-45,8.63982e-46) (1.27141e-44,2.1872e-44) (1.3895e-43,-1.35521e-43) (-1.20625e-42,-7.49e-43) (-3.12136e-42,9.44091e-42) (6.68209e-41,5.86875e-42) (-6.36701e-41,-4.34144e-40) (-2.58136e-39,1.0671e-39) (1.06604e-38,1.35673e-38) (5.70173e-38,-8.51382e-38) (-5.62667e-37,-1.28949e-37) (5.90699e-37,2.98155e-36) (1.14835e-35,-9.21274e-36) (-6.05086e-35,-2.23609e-35) (6.12525e-35,2.44524e-34) (5.33987e-34,-6.83135e-34) (-2.55742e-33,1.79836e-34) (4.80578e-33,4.01593e-33) (-1.84816e-33,-1.20346e-32) (-1.01721e-32,1.60468e-32) (2.42046e-32,-8.97513e-33) (-3.03928e-32,1.84461e-33) (2.95133e-32,-1.42145e-32) (-1.76388e-32,4.18217e-32) (-1.70893e-32,-5.10949e-32) (5.00439e-32,1.65661e-32) (-3.10559e-32,3.30823e-32) (-2.00622e-32,-3.70524e-32) (3.10717e-32,-9.83207e-33) (3.19874e-33,3.44578e-32) (-2.76093e-32,6.03845e-33) (-6.68892e-33,-2.47829e-32) (2.43836e-32,-1.35017e-32) (1.88857e-32,2.82164e-33) (-4.03553e-33,6.98451e-33) (-1.01601e-32,6.22202e-33) (-3.01839e-33,3.15614e-33) (1.45195e-33,1.96389e-35) (1.11408e-33,-8.66726e-34) (1.1143e-34,-3.78565e-34) (-1.23818e-34,1.30669e-35) (-5.43872e-35,6.23153e-35) (-1.05149e-35,1.90217e-35) (-4.81006e-36,-1.73061e-37) (-3.90907e-36,-7.05856e-37) (-1.67008e-36,5.96207e-37) (-2.88783e-37,4.97828e-37) (4.31615e-38,1.4858e-37) (3.32499e-38,1.44245e-38) (6.54256e-39,-3.77608e-39) (9.52981e-41,-1.41954e-39) (-2.00374e-40,-1.42073e-40) (-3.55546e-41,1.66099e-41) (-3.07166e-43,5.82533e-42) (7.04498e-43,4.01322e-43) (8.67729e-44,-6.07429e-44) (-2.47857e-45,-1.28376e-44) (-1.50217e-45,-3.15374e-46) (-9.35942e-47,1.44078e-46) 
  (3.37337e-51,-9.52646e-51) (-1.01735e-49,-1.23238e-50) (1.08952e-49,9.85017e-49) (8.61808e-48,-3.11434e-48) (-4.48373e-47,-6.73097e-47) (-4.58906e-46,5.02423e-46) (4.79387e-45,2.6042e-45) (1.06615e-44,-4.0341e-44) (-3.05317e-43,-7.5052e-45) (4.35171e-43,2.10654e-42) (1.33358e-41,-6.12748e-42) (-6.02339e-41,-7.66507e-41) (-3.80142e-40,5.0258e-40) (3.69016e-39,1.36867e-39) (4.12355e-40,-2.34701e-38) (-1.229e-37,4.78671e-38) (5.01344e-37,4.71953e-37) (8.25405e-37,-3.18538e-36) (-1.35245e-35,4.26175e-36) (4.32999e-35,3.29298e-35) (-4.89532e-36,-1.83106e-34) (-3.7762e-34,3.6805e-34) (1.24857e-33,-1.2712e-35) (-1.77581e-33,-1.55762e-33) (4.56845e-34,3.62572e-33) (2.34964e-33,-4.36387e-33) (-3.65157e-33,4.29142e-33) (1.27274e-33,-5.97702e-33) (4.18082e-33,7.57714e-33) (-9.33018e-33,-3.2686e-33) (7.72412e-33,-5.52971e-33) (1.86019e-33,8.08055e-33) (-7.6711e-33,-8.37594e-34) (1.49562e-33,-5.99571e-33) (5.50813e-33,3.07485e-33) (-1.91527e-33,5.11342e-33) (-4.5753e-33,-1.39028e-33) (7.15793e-34,-4.9527e-33) (2.89904e-33,-2.71287e-33) (6.89037e-34,9.77408e-34) (-4.44195e-34,2.10775e-33) (-1.1979e-35,9.60881e-34) (1.95784e-34,-1.00404e-34) (4.66389e-35,-2.56482e-34) (-3.21866e-35,-7.83284e-35) (-1.61622e-35,1.30185e-35) (5.00383e-37,1.55875e-35) (1.3327e-36,4.53608e-36) (-4.92774e-37,8.39421e-37) (-5.68157e-37,4.80698e-37) (-1.34949e-37,3.19706e-37) (3.15665e-38,1.11351e-37) (2.7712e-38,1.5314e-38) (7.03358e-39,-2.64555e-39) (4.53636e-40,-1.51784e-39) (-1.89141e-40,-2.34584e-40) (-5.2101e-41,6.20489e-42) (-3.34838e-42,7.75633e-42) (7.81057e-43,9.95434e-43) (1.73857e-43,-3.38716e-44) (5.92568e-45,-2.25284e-44) (-2.2414e-45,-1.82873e-45) (-3.02409e-46,1.58165e-46) (4.07935e-48,3.81226e-47) 
  (-4.70735e-52,-2.18274e-51) (-2.04358e-50,9.44392e-51) (1.33238e-49,1.70449e-49) (1.2374e-48,-1.55535e-48) (-1.58154e-47,-7.33043e-48) (-2.83634e-47,1.43077e-46) (1.1642e-45,-4.68168e-47) (-2.38612e-45,-8.58128e-45) (-5.75638e-44,3.11812e-44) (3.06487e-43,3.50571e-43) (1.889e-42,-2.61269e-42) (-2.01878e-41,-8.13241e-42) (-1.56266e-41,1.41694e-40) (8.78096e-40,-1.81664e-40) (-2.86507e-39,-4.51706e-39) (-1.67024e-38,2.47739e-38) (1.53052e-37,1.95692e-38) (-2.78869e-37,-6.70962e-37) (-1.74148e-36,2.53761e-36) (1.15811e-35,-3.33756e-37) (-2.51487e-35,-2.86967e-35) (-1.01715e-35,1.06399e-34) (1.85542e-34,-1.60867e-34) (-4.53634e-34,-1.13749e-35) (5.0983e-34,4.77661e-34) (-2.22424e-34,-9.12389e-34) (1.19643e-34,1.01608e-33) (-7.44228e-34,-8.63015e-34) (1.60606e-33,2.69946e-34) (-1.49603e-33,9.77299e-34) (6.28697e-37,-1.69548e-33) (1.41436e-33,5.38595e-34) (-9.08589e-34,1.05949e-33) (-8.13342e-34,-8.48443e-34) (1.01123e-33,-5.13289e-34) (6.11944e-34,8.46509e-34) (-6.76955e-34,5.87298e-34) (-6.25871e-34,-6.16004e-34) (-5.25586e-35,-7.94098e-34) (1.87898e-34,-6.58589e-35) (2.15806e-34,3.07074e-34) (1.37515e-34,1.46819e-34) (2.48118e-35,-2.64771e-35) (-2.4091e-35,-4.00901e-35) (-1.5583e-35,-8.22241e-36) (-1.33807e-36,3.25919e-36) (2.00224e-36,2.04705e-36) (8.71954e-37,4.77032e-37) (1.01267e-37,1.82627e-37) (3.88392e-39,1.38547e-37) (2.83697e-38,6.08763e-38) (2.03416e-38,1.07977e-38) (6.16237e-39,-1.78518e-39) (6.56016e-40,-1.39704e-39) (-1.48833e-40,-2.93581e-40) (-6.25915e-41,-9.07835e-42) (-7.27854e-42,8.39184e-42) (5.68868e-43,1.71058e-42) (2.67367e-43,5.00979e-44) (2.36944e-44,-3.01599e-44) (-2.19898e-45,-4.57728e-45) (-6.34403e-46,8.58902e-48) (-2.91572e-47,6.93534e-47) (6.03451e-48,5.96493e-48) 
  (-3.36446e-52,-3.52583e-52) (-2.71082e-51,4.06335e-51) (4.36776e-50,1.63803e-50) (5.35198e-50,-4.22529e-49) (-3.6931e-48,3.99602e-49) (1.03211e-47,2.91849e-47) (2.0819e-46,-1.32813e-46) (-1.345e-45,-1.33247e-45) (-7.48957e-45,1.18678e-44) (9.52761e-44,3.41145e-44) (8.0038e-44,-7.07808e-43) (-4.83039e-42,6.99555e-43) (1.36535e-41,2.92467e-41) (1.4566e-40,-1.4226e-40) (-1.10879e-39,-4.85401e-40) (1.46575e-40,6.70198e-39) (2.98669e-38,-1.66341e-38) (-1.37235e-37,-7.9267e-38) (4.41599e-38,6.58082e-37) (1.84481e-36,-1.5897e-36) (-7.74283e-36,-1.21922e-36) (1.21925e-35,1.75359e-35) (7.36006e-36,-4.71125e-35) (-6.78903e-35,5.34791e-35) (1.32459e-34,7.41258e-36) (-1.45917e-34,-9.70886e-35) (1.49258e-34,1.04937e-34) (-2.12263e-34,1.41467e-35) (2.24851e-34,-2.0161e-34) (-2.23994e-35,3.17602e-34) (-2.45509e-34,-1.73025e-34) (2.25018e-34,-1.58966e-34) (6.63836e-35,2.40833e-34) (-2.18985e-34,4.18511e-35) (2.22289e-35,-2.00667e-34) (1.971e-34,-5.85202e-36) (2.43424e-35,1.66748e-34) (-1.48868e-34,2.70963e-35) (-1.24617e-34,-9.06779e-35) (-2.20873e-36,-4.14751e-35) (6.22804e-35,8.04433e-36) (4.03227e-35,1.76717e-36) (3.08064e-36,-6.61863e-36) (-7.7329e-36,-2.5796e-36) (-3.47043e-36,7.81593e-37) (3.81335e-38,6.36738e-37) (5.10491e-37,3.2574e-38) (1.94875e-37,-5.57686e-38) (4.5715e-38,3.89838e-39) (2.08339e-38,1.52e-38) (1.23248e-38,3.6993e-39) (4.30013e-39,-1.4418e-39) (6.15244e-40,-1.13094e-39) (-1.03565e-40,-2.96474e-40) (-6.39032e-41,-2.25501e-41) (-1.08072e-41,7.50193e-42) (6.01959e-44,2.33045e-42) (3.3114e-43,1.89069e-43) (4.98033e-44,-2.96721e-44) (-4.01523e-46,-8.22305e-45) (-1.00395e-45,-4.43147e-46) (-1.04298e-46,9.0303e-47) (4.78221e-48,1.57348e-47) (1.85439e-48,1.73051e-49) 
  (-1.01451e-52,-2.73412e-53) (-4.56851e-53,1.0459e-51) (9.77058e-51,-1.81529e-51) (-3.6185e-50,-8.26563e-50) (-6.28187e-49,4.68353e-49) (4.96079e-48,4.22644e-48) (2.43533e-47,-4.60427e-47) (-3.87341e-46,-1.08252e-46) (-1.792e-46,3.01381e-45) (2.18423e-44,-3.57004e-45) (-6.22491e-44,-1.45574e-43) (-8.54527e-43,6.89051e-43) (6.11608e-42,3.98149e-42) (9.90185e-42,-4.49028e-41) (-2.66708e-40,5.12558e-41) (8.94907e-40,1.18932e-39) (3.05774e-39,-6.83321e-39) (-3.38342e-38,4.57459e-39) (9.40463e-38,1.0312e-37) (8.74841e-38,-4.97522e-37) (-1.36164e-36,8.17002e-37) (4.06678e-36,1.08631e-36) (-4.73438e-36,-7.83083e-36) (-3.45171e-36,1.59661e-35) (1.99424e-35,-1.50668e-35) (-3.17029e-35,5.41546e-36) (3.10442e-35,-7.87796e-36) (-2.17488e-35,3.32464e-35) (-3.09578e-36,-5.50209e-35) (4.23892e-35,3.65737e-35) (-4.9699e-35,1.8187e-35) (-1.00142e-36,-4.99049e-35) (4.2192e-35,1.3768e-35) (-1.63184e-35,3.86485e-35) (-2.78695e-35,-2.24389e-35) (1.98835e-35,-3.08176e-35) (2.86677e-35,1.33765e-35) (-1.02324e-35,2.36776e-35) (-2.80412e-35,6.93597e-36) (-8.90378e-36,-3.6436e-36) (7.56711e-36,-6.58226e-36) (5.77401e-36,-5.23902e-36) (-1.91324e-38,-1.66457e-36) (-1.28937e-36,4.94664e-37) (-4.14508e-37,5.6158e-37) (6.16474e-38,1.09937e-37) (7.0347e-38,-5.41935e-38) (1.98773e-38,-3.49439e-38) (6.68238e-39,-7.48713e-39) (4.61235e-39,-1.40585e-39) (2.07109e-39,-1.29713e-39) (3.69109e-40,-8.03632e-40) (-7.47204e-41,-2.44744e-40) (-5.68313e-41,-2.79064e-41) (-1.25903e-41,5.71234e-42) (-5.66742e-43,2.6524e-42) (3.37144e-43,3.48627e-43) (7.81318e-44,-1.7024e-44) (3.72098e-45,-1.16701e-44) (-1.21429e-45,-1.26303e-45) (-2.25056e-46,6.80858e-47) (-4.59065e-48,2.93878e-47) (2.98084e-48,1.95543e-48) (3.35695e-49,-2.2745e-49) 
  (-2.15245e-53,6.12504e-54) (1.05287e-52,1.95114e-52) (1.57545e-51,-1.37801e-51) (-1.53032e-50,-1.1125e-50) (-6.50173e-50,1.50464e-49) (1.33965e-48,2.60547e-49) (-2.01238e-49,-1.09711e-47) (-8.3529e-47,1.92381e-47) (2.78261e-46,5.91703e-46) (3.82346e-45,-3.02536e-45) (-2.82971e-44,-2.12041e-44) (-8.40777e-44,2.32285e-43) (1.64388e-42,1.50463e-44) (-3.76102e-42,-9.60019e-42) (-4.20013e-41,4.33568e-41) (3.12719e-40,9.50705e-41) (-3.64565e-40,-1.57829e-39) (-5.07639e-39,5.19681e-39) (2.88093e-38,4.51352e-39) (-5.08478e-38,-9.00496e-38) (-1.03639e-37,2.99921e-37) (7.40701e-37,-3.48735e-37) (-1.64299e-36,-5.64703e-37) (1.40903e-36,2.72311e-36) (9.88775e-37,-4.55868e-36) (-3.42963e-36,4.67093e-36) (2.35908e-36,-5.02886e-36) (2.47436e-36,6.97828e-36) (-8.05425e-36,-5.73059e-36) (9.48482e-36,-2.1844e-36) (-2.29148e-36,9.00452e-36) (-7.5211e-36,-4.9076e-36) (6.1102e-36,-4.93719e-36) (4.22338e-36,6.55659e-36) (-5.99157e-36,2.09345e-36) (-2.56578e-36,-6.20908e-36) (5.05845e-36,-3.03271e-36) (2.49138e-36,3.62547e-36) (-2.31534e-36,4.70839e-36) (-1.79065e-36,1.25923e-36) (-2.1707e-38,-1.51415e-36) (7.04166e-38,-1.45188e-36) (-2.11126e-37,-3.16345e-37) (-1.1802e-37,1.95075e-37) (1.06614e-38,1.32864e-37) (2.24544e-38,1.39191e-38) (3.14211e-39,-1.46259e-38) (-1.94844e-39,-7.51858e-39) (-3.41177e-40,-2.12704e-39) (3.03633e-40,-8.58324e-40) (6.97212e-41,-4.55416e-40) (-6.5194e-41,-1.5788e-40) (-4.47903e-41,-2.30802e-41) (-1.19862e-41,4.04063e-42) (-1.02868e-42,2.59951e-42) (2.87672e-43,4.73786e-43) (9.98664e-44,5.6739e-45) (9.66799e-45,-1.35273e-44) (-1.04279e-45,-2.34478e-45) (-3.68349e-46,-3.17202e-47) (-2.67621e-47,4.21809e-47) (3.32089e-48,5.42325e-48) (7.61228e-49,-8.92509e-50) (2.45984e-50,-8.40513e-50) 
  (-3.24333e-54,3.41571e-54) (3.96915e-53,2.40752e-53) (1.39937e-52,-4.13261e-52) (-3.90981e-51,-4.3152e-52) (3.4803e-51,3.39172e-50) (2.71803e-49,-8.68034e-50) (-1.13717e-48,-2.02055e-48) (-1.38422e-47,1.21145e-47) (1.15181e-46,8.44135e-47) (4.0931e-46,-1.00074e-45) (-7.8701e-45,-8.66657e-46) (1.15036e-44,5.42776e-44) (3.10048e-43,-1.98579e-43) (-1.89548e-42,-1.28937e-42) (-1.98404e-42,1.31311e-41) (6.68505e-41,-2.38075e-41) (-2.66917e-40,-2.20638e-40) (-1.62837e-40,1.51811e-39) (5.20981e-39,-3.0091e-39) (-1.95066e-38,-7.48737e-39) (2.23591e-38,5.84325e-38) (6.57355e-38,-1.42837e-37) (-3.05452e-37,1.15794e-37) (5.26148e-37,2.2347e-37) (-4.16295e-37,-7.5362e-37) (1.5041e-37,1.01282e-36) (-4.32033e-37,-8.54014e-37) (1.30355e-36,4.28268e-37) (-1.67397e-36,4.81106e-37) (6.47462e-37,-1.54678e-36) (1.08006e-36,1.21723e-36) (-1.48014e-36,6.12055e-37) (-1.537e-37,-1.38198e-36) (1.42786e-36,4.90587e-38) (-2.40526e-37,1.10599e-36) (-1.18502e-36,-2.58342e-37) (7.08924e-38,-1.08484e-36) (7.58987e-37,-4.85828e-38) (3.74924e-37,8.44858e-37) (-1.32238e-38,4.73826e-37) (-1.70929e-37,-1.27172e-37) (-1.7675e-37,-1.93158e-37) (-7.89079e-38,-2.67129e-38) (2.85948e-39,3.68415e-38) (1.77151e-38,1.73664e-38) (5.61468e-39,-7.98636e-41) (-1.09822e-39,-2.18206e-39) (-1.24701e-39,-7.65394e-40) (-3.84319e-40,-2.36814e-40) (-9.77734e-41,-1.43987e-40) (-5.66628e-41,-6.52029e-41) (-3.07024e-41,-1.12566e-41) (-9.30987e-42,3.15925e-42) (-1.11326e-42,2.24355e-42) (2.1521e-43,5.17371e-43) (1.08339e-43,2.95406e-44) (1.57602e-44,-1.30399e-44) (-4.02392e-46,-3.40458e-45) (-4.86166e-46,-2.1881e-46) (-6.2261e-47,4.59218e-47) (1.55684e-48,1.0409e-47) (1.28211e-48,4.17468e-49) (1.1196e-49,-1.19067e-49) (-7.44434e-51,-1.72245e-50) 
  (-2.26888e-55,9.53673e-55) (9.61802e-54,2.31911e-55) (-1.68477e-53,-8.85907e-53) (-7.50127e-52,3.13774e-52) (3.99331e-51,5.84499e-51) (4.17351e-50,-4.28563e-50) (-4.14932e-49,-2.66984e-49) (-1.40792e-48,3.72745e-48) (3.11842e-47,4.04984e-48) (-3.22223e-47,-2.38688e-46) (-1.60737e-45,7.47211e-46) (8.69441e-45,8.85118e-45) (3.27733e-44,-7.50019e-44) (-5.04848e-43,5.86522e-45) (1.32691e-42,2.56764e-42) (8.41478e-42,-1.2693e-41) (-7.31067e-41,-2.41414e-42) (1.6935e-40,2.67936e-40) (4.37537e-40,-1.14501e-39) (-3.94804e-39,1.33248e-39) (1.0642e-38,5.91329e-39) (-7.85118e-39,-2.87923e-38) (-3.01002e-38,5.29302e-38) (1.01334e-37,-3.05466e-38) (-1.47942e-37,-5.22147e-38) (1.4333e-37,1.04309e-37) (-1.62522e-37,-2.84663e-38) (2.09737e-37,-1.39482e-37) (-1.14118e-37,2.78953e-37) (-1.52841e-37,-2.4301e-37) (2.81918e-37,-3.74244e-38) (-5.87711e-38,2.76694e-37) (-2.21743e-37,-1.0838e-37) (1.54878e-37,-2.05816e-37) (1.46836e-37,1.40659e-37) (-1.57915e-37,1.47469e-37) (-1.5369e-37,-1.24051e-37) (6.02856e-38,-1.20403e-37) (1.52226e-37,4.23122e-38) (7.42383e-38,6.34595e-38) (-2.55591e-38,1.02523e-38) (-4.55166e-38,-1.65516e-39) (-1.6198e-38,6.35799e-39) (3.61621e-39,4.7595e-39) (4.49665e-39,2.86501e-40) (9.48171e-40,-6.97134e-40) (-3.46195e-40,-1.72992e-40) (-2.62868e-40,5.6606e-41) (-8.84564e-41,2.61316e-41) (-3.36198e-41,-1.47224e-42) (-1.61351e-41,3.10384e-43) (-5.50207e-42,2.87857e-42) (-8.03463e-43,1.72326e-42) (1.58371e-43,4.65385e-43) (1.02444e-43,4.36211e-44) (1.98432e-44,-1.07247e-44) (5.33518e-46,-4.11351e-45) (-5.30464e-46,-4.58279e-46) (-1.04652e-46,3.33878e-47) (-3.37306e-48,1.56975e-47) (1.67313e-48,1.42738e-48) (2.61844e-49,-1.08842e-49) (1.83377e-51,-3.45229e-50) (-3.5598e-51,-1.79975e-51) 
  (5.62664e-56,1.93969e-55) (1.74879e-54,-9.22413e-55) (-1.17861e-53,-1.43007e-53) (-1.05767e-52,1.30208e-52) (1.30247e-51,6.89652e-52) (3.63444e-51,-1.21002e-50) (-1.05654e-49,-9.3932e-51) (1.15484e-49,8.63874e-49) (6.46454e-48,-2.60367e-48) (-3.32946e-47,-4.21833e-47) (-2.16438e-46,3.31225e-46) (2.69295e-45,5.8982e-46) (-3.3504e-45,-1.77233e-44) (-8.90224e-44,6.47223e-44) (5.57324e-43,2.76273e-43) (-2.04019e-43,-3.22359e-42) (-1.23438e-41,8.98064e-42) (6.14252e-41,2.12674e-41) (-7.74589e-41,-2.34139e-40) (-4.30185e-40,6.98465e-40) (2.29685e-39,-4.42922e-40) (-4.59453e-39,-3.20551e-39) (1.939e-39,1.1093e-38) (1.06485e-38,-1.62725e-38) (-2.59953e-38,1.08776e-38) (2.95637e-38,-5.38726e-39) (-2.05229e-38,2.00173e-38) (3.98745e-39,-4.54704e-38) (2.55122e-38,4.44285e-38) (-4.8939e-38,-2.0877e-39) (2.20741e-38,-4.43776e-38) (3.41102e-38,3.58116e-38) (-3.74884e-38,2.29753e-38) (-1.41194e-38,-4.34629e-38) (3.56034e-38,-9.14776e-39) (5.65884e-39,3.7627e-38) (-3.39972e-38,9.5062e-39) (-1.32165e-38,-2.05539e-38) (2.12913e-38,-1.52985e-38) (1.89964e-38,-3.11464e-39) (2.47024e-40,3.44058e-39) (-5.53063e-39,5.26901e-39) (-1.57561e-39,3.10104e-39) (9.14974e-40,3.85027e-40) (6.40472e-40,-4.7894e-40) (6.71204e-41,-2.3098e-40) (-5.94772e-41,7.34841e-42) (-2.72414e-41,3.97706e-41) (-8.13599e-42,1.64845e-41) (-4.20277e-42,5.02944e-42) (-1.87137e-42,2.35676e-42) (-2.89315e-43,1.13419e-42) (1.33743e-43,3.39203e-43) (8.6122e-44,4.16549e-44) (2.04159e-44,-8.0273e-45) (1.37384e-45,-4.27737e-45) (-4.87559e-46,-6.76819e-46) (-1.42101e-46,4.34947e-48) (-1.13079e-47,1.93936e-47) (1.62564e-48,2.87765e-48) (4.55806e-49,-5.43319e-51) (2.65769e-50,-5.28479e-50) (-4.39418e-51,-5.77237e-51) (-8.19425e-52,1.90792e-52) 
  (2.92017e-56,2.91654e-56) (2.24664e-55,-3.35868e-55) (-3.50962e-54,-1.46087e-54) (-7.00649e-54,3.39968e-53) (3.09189e-52,3.95338e-54) (-4.93434e-52,-2.65234e-51) (-2.12691e-50,8.90821e-51) (1.14031e-49,1.54732e-49) (9.55381e-49,-1.22025e-48) (-1.1222e-47,-4.17377e-48) (-8.88322e-49,8.78497e-47) (5.65797e-46,-2.21709e-46) (-2.80858e-45,-2.7585e-45) (-7.41881e-45,2.25493e-44) (1.30241e-43,-2.36163e-44) (-4.44738e-43,-5.1051e-43) (-8.57875e-43,3.02852e-42) (1.24001e-41,-4.43501e-42) (-4.13962e-41,-2.62257e-41) (2.25743e-41,1.57845e-40) (2.80396e-40,-3.44243e-40) (-1.03736e-39,8.74872e-41) (1.57084e-39,1.34443e-39) (-4.3947e-40,-3.51531e-39) (-2.07677e-39,4.52818e-39) (2.66455e-39,-4.21609e-39) (7.89723e-40,4.98293e-39) (-5.85481e-39,-5.65748e-39) (8.49138e-39,1.11069e-39) (-4.98638e-39,6.69781e-39) (-4.23566e-39,-7.49002e-39) (8.45244e-39,-1.39296e-39) (-1.70941e-40,7.8494e-39) (-7.63999e-39,-2.32333e-39) (2.05843e-39,-6.33754e-39) (5.9797e-39,2.88059e-39) (-2.11677e-39,5.8314e-39) (-4.50559e-39,7.04464e-41) (1.48372e-40,-4.22537e-39) (1.90902e-39,-3.10793e-39) (5.84644e-40,-1.40735e-41) (-8.56294e-42,1.23058e-39) (1.80032e-40,6.43455e-40) (1.7337e-40,-1.70991e-41) (3.19257e-41,-1.35226e-40) (-1.83145e-41,-4.41683e-41) (-7.49265e-42,5.501e-42) (1.28026e-42,8.32813e-42) (1.2467e-42,3.35265e-42) (2.6284e-43,1.25142e-42) (1.18714e-43,5.48201e-43) (1.22796e-43,1.81596e-43) (6.44399e-44,2.56537e-44) (1.73713e-44,-6.25336e-45) (1.73132e-45,-3.92099e-45) (-3.91259e-46,-7.9649e-46) (-1.63357e-46,-3.15191e-47) (-2.0407e-47,2.00365e-47) (9.42375e-49,4.45246e-48) (6.38831e-49,2.17692e-49) (6.96958e-50,-6.2666e-50) (-2.99423e-51,-1.18702e-50) (-1.4758e-51,-3.21145e-52) (-1.05589e-52,1.40918e-52) 
  (8.02797e-57,2.44263e-57) (8.94165e-57,-8.19879e-56) (-7.80076e-55,6.12917e-56) (1.89335e-54,6.99026e-54) (5.89487e-53,-2.88932e-53) (-3.58094e-52,-4.60479e-52) (-3.18801e-51,3.93281e-51) (3.8872e-50,1.74424e-50) (4.38219e-50,-3.41828e-49) (-2.60176e-48,5.35645e-49) (1.04464e-47,1.63084e-47) (7.48165e-47,-1.09646e-46) (-8.39414e-46,-1.36271e-46) (1.5593e-45,4.81779e-45) (1.89073e-44,-2.04409e-44) (-1.37566e-43,-2.73657e-44) (2.4572e-43,5.9243e-43) (1.37306e-42,-2.25018e-42) (-9.54429e-42,1.18585e-42) (2.27221e-41,2.05109e-41) (-9.95213e-43,-8.32919e-41) (-1.36861e-40,1.34185e-40) (3.76936e-40,6.46207e-42) (-4.73434e-40,-4.29275e-40) (2.75136e-40,8.2072e-40) (-2.27599e-40,-7.78491e-40) (8.05891e-40,3.994e-40) (-1.41637e-39,1.66882e-40) (9.80282e-40,-1.01423e-39) (4.71212e-40,1.34386e-39) (-1.48111e-39,-1.20701e-40) (6.14209e-40,-1.33783e-39) (1.15508e-39,7.93038e-40) (-1.07813e-39,8.56272e-40) (-7.56926e-40,-9.38198e-40) (9.93e-40,-5.78314e-40) (6.08442e-40,8.83152e-40) (-4.47356e-40,7.03308e-40) (-5.22478e-40,-4.10853e-40) (-1.96972e-40,-6.3694e-40) (3.30661e-41,-1.38124e-40) (1.36125e-40,1.31419e-40) (1.05836e-40,6.40871e-41) (2.65917e-41,-1.8604e-41) (-1.03714e-41,-2.12882e-41) (-8.16879e-42,-4.34e-42) (-7.37332e-43,1.32964e-42) (1.12326e-42,8.92002e-43) (6.24225e-43,2.69969e-43) (2.20826e-43,1.14043e-43) (9.31506e-44,4.75135e-44) (4.04963e-44,5.17274e-45) (1.18353e-44,-5.59993e-45) (1.45861e-45,-3.21932e-45) (-2.98687e-46,-7.7508e-46) (-1.63678e-46,-5.86152e-47) (-2.77454e-47,1.77072e-47) (-2.64551e-49,5.701e-48) (7.43156e-49,5.34341e-49) (1.25828e-49,-5.34956e-50) (2.20975e-51,-1.8991e-50) (-2.06243e-51,-1.43683e-51) (-2.74728e-52,1.47863e-52) (2.12236e-54,3.65107e-53) 
  (1.67812e-57,-3.0258e-58) (-5.91403e-57,-1.58345e-56) (-1.39452e-55,8.34766e-56) (1.0159e-54,1.14468e-54) (8.50578e-54,-1.12845e-53) (-1.16201e-52,-5.26563e-53) (-1.9634e-52,1.1016e-51) (9.40444e-51,-9.98086e-52) (-3.13281e-50,-6.96747e-50) (-4.18708e-49,4.09328e-49) (3.88035e-48,1.6915e-48) (-2.38603e-49,-2.87083e-47) (-1.62728e-46,8.09542e-47) (8.6875e-46,6.21555e-46) (5.58641e-46,-5.76335e-45) (-2.5665e-44,1.28856e-44) (1.13004e-43,6.25223e-44) (-6.95755e-44,-5.16674e-43) (-1.28122e-42,1.35471e-42) (5.80083e-42,2.31665e-43) (-1.00276e-41,-1.17635e-41) (-3.68075e-42,3.47975e-41) (5.32593e-41,-4.26893e-41) (-1.13989e-40,-2.28054e-42) (1.30635e-40,6.87789e-41) (-1.18689e-40,-5.19423e-41) (1.43187e-40,-7.51046e-41) (-1.32178e-40,2.0619e-40) (-4.11304e-41,-2.26028e-40) (2.35057e-40,6.14961e-41) (-1.6003e-40,1.98518e-40) (-1.31711e-40,-2.14223e-40) (2.31241e-40,-9.22768e-41) (1.73152e-41,2.34196e-40) (-2.15817e-40,1.91834e-41) (1.26812e-41,-1.97388e-40) (1.82641e-40,2.09773e-42) (5.91211e-41,1.41023e-40) (-9.77424e-41,3.13591e-41) (-1.07448e-40,-4.83676e-41) (-2.4975e-41,-2.36357e-41) (2.74096e-41,-1.48191e-42) (2.16125e-41,-4.74668e-42) (2.45135e-42,-5.7602e-42) (-3.58168e-42,-1.71558e-42) (-1.70651e-42,3.61658e-43) (-2.86842e-44,2.7448e-43) (2.36803e-43,-1.62433e-44) (1.16836e-43,-4.83582e-44) (4.42146e-44,-1.84504e-44) (1.78555e-44,-7.82888e-45) (5.65711e-45,-5.0247e-45) (7.33983e-46,-2.34175e-45) (-2.47913e-46,-6.23861e-46) (-1.46071e-46,-6.45359e-47) (-3.07218e-47,1.40667e-47) (-1.54412e-48,6.27256e-48) (7.31705e-49,8.61002e-49) (1.8138e-49,-2.1483e-50) (1.16087e-50,-2.49112e-50) (-2.21369e-51,-3.17406e-51) (-5.09064e-52,5.56554e-53) (-2.29399e-53,5.96964e-53) (5.2005e-54,5.45717e-54) 
  (2.80082e-58,-2.0713e-58) (-2.5377e-57,-2.40981e-57) (-1.86799e-56,2.86859e-56) (3.04511e-55,1.22774e-55) (5.19815e-55,-3.03685e-54) (-2.80578e-53,1.99361e-54) (8.32989e-53,2.33566e-52) (1.67099e-51,-1.2632e-51) (-1.40333e-50,-9.30467e-51) (-2.72874e-50,1.25094e-49) (9.00232e-49,-1.71369e-49) (-3.58575e-48,-4.99041e-48) (-1.77507e-47,3.4077e-47) (2.22761e-46,-4.68534e-48) (-6.29818e-46,-1.01009e-45) (-2.47729e-45,5.25753e-45) (2.53327e-44,-4.33956e-45) (-7.43246e-44,-6.96889e-44) (-2.38821e-44,3.56358e-43) (8.63655e-43,-6.62027e-43) (-2.79702e-42,-4.87578e-43) (3.49311e-42,5.28971e-42) (2.42636e-42,-1.20246e-41) (-1.53207e-41,1.29936e-41) (2.36683e-41,-7.00752e-42) (-1.80093e-41,9.66334e-42) (4.62947e-42,-2.87223e-41) (1.27212e-41,3.91667e-41) (-3.38913e-41,-1.53229e-41) (3.11467e-41,-2.72892e-41) (1.26224e-41,4.15677e-41) (-4.27756e-41,-1.44008e-42) (9.53827e-42,-4.2851e-41) (3.45905e-41,1.96032e-41) (-1.89027e-41,3.36031e-41) (-2.68974e-41,-2.06147e-41) (1.78314e-41,-2.50206e-41) (2.68753e-41,6.31617e-42) (-3.71337e-42,1.53883e-41) (-1.83669e-41,8.31702e-42) (-7.53771e-42,1.31504e-42) (2.29055e-42,-2.87815e-42) (2.12455e-42,-3.18017e-42) (-2.48675e-43,-1.18705e-42) (-6.44162e-43,1.35526e-43) (-1.97183e-43,2.53656e-43) (1.8626e-44,5.16495e-44) (2.65765e-44,-2.72636e-44) (8.57916e-45,-2.13402e-44) (2.84223e-45,-8.6768e-45) (9.89494e-46,-3.49476e-45) (-1.67619e-47,-1.39636e-45) (-2.29188e-46,-3.95268e-46) (-1.17284e-46,-4.75399e-47) (-2.83541e-47,1.1137e-47) (-2.32658e-48,6.08587e-48) (6.28059e-49,1.08986e-48) (2.20548e-49,2.50356e-50) (2.35514e-50,-2.74452e-50) (-1.61447e-51,-5.23869e-51) (-7.55916e-52,-1.80775e-52) (-6.99889e-53,7.62906e-53) (4.40503e-54,1.22408e-53) (1.5338e-54,1.60213e-55) 
  (3.37602e-59,-6.35948e-59) (-7.00036e-58,-2.26187e-58) (-8.9625e-58,7.27325e-57) (7.11718e-56,-6.12359e-57) (-2.12837e-55,-6.43818e-55) (-5.20025e-54,3.42265e-54) (4.21745e-53,3.51255e-53) (1.66253e-52,-4.30645e-52) (-3.68271e-51,-4.07593e-53) (1.02119e-50,2.5791e-50) (1.37454e-49,-1.40259e-49) (-1.23269e-48,-4.16953e-49) (1.23569e-48,7.93787e-48) (3.60804e-47,-2.84593e-47) (-2.26824e-46,-8.41289e-47) (2.62769e-46,1.13262e-45) (3.34768e-45,-3.78855e-45) (-1.96327e-44,-1.33411e-45) (3.95147e-44,5.48557e-44) (4.47404e-44,-1.96668e-43) (-4.48788e-43,2.55818e-43) (1.08977e-42,3.35004e-43) (-1.05046e-42,-1.91805e-42) (-4.76932e-43,3.45871e-42) (1.93632e-42,-3.54612e-42) (-4.42102e-43,3.1856e-42) (-3.55125e-42,-3.79874e-42) (6.31763e-42,2.44186e-42) (-5.10812e-42,3.19589e-42) (-8.4277e-43,-6.98287e-42) (7.0148e-42,2.18586e-42) (-4.19939e-42,5.93627e-42) (-5.19467e-42,-5.62893e-42) (5.96873e-42,-3.05833e-42) (2.93929e-42,6.10532e-42) (-5.47527e-42,1.85964e-42) (-1.76854e-42,-4.80698e-42) (3.74374e-42,-3.13549e-42) (1.85232e-42,1.68415e-42) (-9.68617e-43,3.19786e-42) (-7.85669e-43,1.37473e-42) (-9.80106e-44,-4.24688e-43) (-1.14389e-43,-6.28163e-43) (-1.74898e-43,-1.51411e-43) (-7.20854e-44,8.1046e-44) (2.40773e-45,5.78494e-44) (8.67031e-45,7.25033e-45) (3.3673e-46,-5.88506e-45) (-1.6338e-45,-3.75353e-45) (-8.69902e-46,-1.47984e-45) (-3.81653e-46,-5.56885e-46) (-1.96366e-46,-1.65425e-46) (-8.26403e-47,-1.78236e-47) (-2.15678e-47,9.78834e-48) (-2.26115e-48,5.30548e-48) (5.01676e-49,1.1413e-48) (2.33514e-49,6.74122e-50) (3.46289e-50,-2.59428e-50) (-2.62814e-52,-7.10142e-51) (-9.33766e-52,-5.52752e-52) (-1.36358e-52,7.35323e-53) (-4.28131e-55,2.07683e-53) (2.29107e-54,1.28422e-54) (2.5783e-55,-1.77706e-55) 
  (7.29731e-61,-1.51161e-59) (-1.55936e-58,2.12567e-59) (5.31072e-58,1.50162e-57) (1.32391e-56,-8.44698e-57) (-1.09986e-55,-1.01906e-55) (-6.13828e-55,1.2328e-54) (1.19642e-53,1.76457e-54) (-1.99682e-53,-9.90011e-53) (-6.7051e-52,4.33397e-52) (4.93332e-51,3.32652e-51) (6.65968e-51,-4.11069e-50) (-2.60286e-49,8.09514e-50) (1.18491e-48,1.16416e-48) (2.33499e-48,-9.07607e-48) (-4.63466e-47,1.46646e-47) (1.8e-46,1.43108e-46) (4.33629e-47,-9.82121e-46) (-3.05983e-45,2.17906e-45) (1.22399e-44,3.19341e-45) (-1.66946e-44,-3.30018e-44) (-3.31259e-44,8.70849e-44) (1.88223e-43,-7.77103e-44) (-3.60973e-43,-1.37804e-43) (3.37709e-43,4.93294e-43) (-1.88348e-43,-6.18501e-43) (3.80511e-43,3.43065e-43) (-9.14889e-43,7.11853e-44) (9.41563e-43,-5.47505e-43) (-1.40107e-44,9.83335e-43) (-1.05127e-42,-5.52001e-43) (9.64864e-43,-7.69807e-43) (4.50865e-43,1.14941e-42) (-1.30836e-42,1.75316e-43) (1.15586e-43,-1.12512e-42) (1.15821e-42,1.95471e-43) (-2.55489e-43,9.48744e-43) (-8.25765e-43,-2.00141e-43) (-3.78457e-44,-8.43486e-43) (3.9076e-43,-1.45204e-43) (2.86673e-43,4.53047e-43) (1.01454e-43,2.92323e-43) (-4.02529e-44,-1.06244e-44) (-8.36718e-44,-5.96365e-44) (-4.30045e-44,-1.38316e-45) (-1.89994e-45,1.77851e-44) (6.92044e-45,7.5311e-45) (2.29649e-45,2.38695e-46) (-5.20253e-46,-7.04025e-46) (-6.64681e-46,-2.57664e-46) (-3.116e-46,-6.32349e-47) (-1.24358e-46,-1.23836e-47) (-4.64379e-47,7.47816e-48) (-1.26229e-47,9.08374e-48) (-1.4267e-48,4.16454e-48) (4.16166e-49,1.00075e-48) (2.20363e-49,8.6569e-50) (4.11504e-50,-2.18822e-50) (1.40944e-51,-8.25135e-51) (-9.80212e-52,-9.79683e-52) (-2.08709e-52,4.34452e-53) (-1.03563e-53,2.88457e-53) (2.6754e-54,3.15512e-54) (5.15216e-55,-1.07513e-55) (1.6082e-56,-6.10334e-56) 
  (-1.24333e-60,-2.99299e-60) (-2.83805e-59,1.91003e-59) (2.55045e-58,2.39744e-58) (1.67799e-57,-3.03831e-57) (-3.23074e-56,-7.45317e-57) (2.41723e-56,3.02439e-55) (2.42199e-54,-1.06618e-54) (-1.53661e-53,-1.56088e-53) (-6.7184e-53,1.57663e-52) (1.26291e-51,-1.89443e-53) (-3.88272e-51,-7.82557e-51) (-3.35504e-50,4.5431e-50) (3.36729e-49,4.47527e-50) (-7.41559e-49,-1.73838e-48) (-5.44994e-48,7.97369e-48) (4.4967e-47,-8.61013e-50) (-1.12449e-46,-1.5189e-46) (-1.85187e-46,6.84264e-46) (2.1215e-45,-9.88266e-46) (-6.15249e-45,-2.68666e-45) (5.31809e-45,1.57997e-44) (1.69239e-44,-3.19098e-44) (-6.3589e-44,2.29094e-44) (9.81568e-44,2.25895e-44) (-9.02798e-44,-4.5297e-44) (8.09752e-44,-2.19912e-44) (-9.09695e-44,1.30593e-43) (2.32775e-44,-1.697e-43) (1.35808e-43,8.91661e-44) (-1.76276e-43,9.18473e-44) (-1.65315e-44,-2.05507e-43) (2.04983e-43,4.3524e-44) (-1.04085e-43,1.98918e-43) (-1.49149e-43,-1.1957e-43) (1.42128e-43,-1.41721e-43) (1.08967e-43,1.25437e-43) (-1.03057e-43,9.59652e-44) (-1.16669e-43,-8.19321e-44) (9.92058e-45,-7.27056e-44) (8.24319e-44,1.13586e-44) (5.32081e-44,2.23253e-44) (2.16192e-46,4.18384e-45) (-1.56875e-44,2.42923e-45) (-6.08972e-45,4.83128e-45) (1.43194e-45,2.60167e-45) (1.75949e-45,2.27073e-46) (3.96617e-46,-2.33887e-46) (-1.189e-46,-3.39347e-47) (-1.10887e-46,4.94159e-47) (-4.67736e-47,3.42498e-47) (-1.65891e-47,1.59273e-47) (-4.49712e-48,7.31143e-48) (-3.06885e-49,2.82851e-48) (3.81084e-49,7.17896e-49) (1.88074e-49,7.43452e-50) (4.09144e-50,-1.78334e-50) (2.70154e-51,-8.4494e-51) (-8.97132e-52,-1.33373e-51) (-2.68109e-52,-9.10248e-54) (-2.42727e-53,3.37512e-53) (2.28328e-54,5.56857e-54) (8.09568e-55,1.15223e-55) (6.305e-56,-8.35786e-56) (-5.54103e-57,-1.13488e-56) 
  (-5.28288e-61,-4.67769e-61) (-3.64959e-60,6.57659e-60) (7.47386e-59,1.99668e-59) (-8.25813e-60,-7.67319e-58) (-6.95662e-57,2.22479e-57) (3.93948e-56,5.34431e-56) (3.16212e-55,-4.79143e-55) (-4.60586e-54,-9.57275e-55) (7.21586e-54,3.56874e-53) (2.14325e-52,-1.56309e-52) (-1.60525e-51,-8.42347e-52) (2.32529e-53,1.1574e-50) (5.97412e-50,-3.3928e-50) (-3.29132e-49,-1.83698e-49) (1.29108e-49,1.8932e-48) (6.77309e-48,-5.45218e-48) (-3.47996e-47,-8.90685e-48) (5.44141e-47,1.20557e-46) (1.84075e-46,-3.86767e-46) (-1.16095e-45,3.3092e-46) (2.51089e-45,1.56882e-45) (-1.30555e-45,-6.22551e-45) (-5.69649e-45,1.02126e-44) (1.4432e-44,-8.36011e-45) (-1.43793e-44,5.47538e-45) (4.24865e-45,-1.35828e-44) (7.15037e-45,2.6082e-44) (-1.87342e-44,-1.85813e-44) (2.48053e-44,-1.11e-44) (-4.20878e-45,3.26735e-44) (-2.9909e-44,-1.6759e-44) (2.5385e-44,-2.48408e-44) (1.71538e-44,3.35461e-44) (-3.07565e-44,1.01948e-44) (-5.48035e-45,-3.33655e-44) (2.77414e-44,-3.35037e-45) (3.96145e-45,2.30491e-44) (-2.24455e-44,6.97668e-45) (-1.0471e-44,-8.28358e-45) (9.12183e-45,-8.51471e-45) (9.3755e-45,-4.35168e-45) (1.3316e-45,-2.10574e-46) (-1.40317e-45,1.86959e-45) (-2.47334e-46,1.33943e-45) (4.4601e-46,2.21603e-46) (2.55205e-46,-1.62718e-46) (3.26178e-47,-8.3143e-47) (-1.57058e-47,5.00491e-48) (-7.17161e-48,1.88827e-47) (-1.15883e-48,1.03353e-47) (2.1926e-49,4.19397e-48) (4.71733e-49,1.48678e-48) (3.46448e-49,3.84772e-49) (1.44034e-49,3.85669e-50) (3.41099e-50,-1.55195e-50) (3.03142e-51,-7.78398e-51) (-7.53056e-52,-1.49739e-51) (-2.99359e-52,-6.52717e-53) (-3.87622e-53,3.39821e-53) (9.71513e-55,7.98921e-54) (1.0587e-54,5.05652e-55) (1.33611e-55,-8.88692e-56) (-1.5416e-57,-2.06167e-56) (-2.30825e-57,-9.83012e-58) 
  (-1.50299e-61,-3.93561e-62) (-2.80865e-62,1.66263e-60) (1.65704e-59,-4.23349e-60) (-8.725e-59,-1.44754e-58) (-1.04262e-57,1.21127e-57) (1.3441e-56,5.18148e-57) (4.09009e-59,-1.2334e-55) (-9.24164e-55,3.82003e-55) (5.5382e-54,5.28234e-54) (1.73083e-53,-5.23266e-53) (-3.68016e-52,5.52179e-53) (1.40972e-51,1.87548e-51) (5.37598e-51,-1.26489e-50) (-7.34847e-50,1.1304e-50) (2.48163e-49,2.72712e-49) (3.55094e-49,-1.62429e-48) (-6.12701e-48,2.83681e-48) (2.18899e-47,1.07974e-47) (-1.88674e-47,-7.52547e-47) (-1.22382e-46,1.76981e-46) (5.17792e-46,-6.73687e-47) (-8.73958e-46,-6.8693e-46) (4.2297e-46,1.9536e-45) (7.68488e-46,-2.59975e-45) (-7.90303e-46,2.14332e-45) (-1.56573e-45,-1.92777e-45) (4.07877e-45,1.88317e-45) (-3.94083e-45,6.73844e-46) (7.2238e-46,-4.52629e-45) (4.0053e-45,3.6258e-45) (-5.06553e-45,2.57632e-45) (-1.08646e-45,-5.90208e-45) (6.18134e-45,8.827e-46) (-1.41605e-45,5.31641e-45) (-5.04014e-45,-2.48397e-45) (2.14605e-45,-4.1471e-45) (3.57313e-45,1.55397e-45) (-1.3033e-45,3.55493e-45) (-2.31717e-45,7.6864e-46) (-1.74843e-46,-1.79902e-45) (5.4193e-46,-1.70162e-45) (1.43716e-46,-3.52168e-46) (4.1549e-47,3.21115e-46) (1.19847e-46,1.97805e-46) (8.33016e-47,-1.26789e-47) (1.55756e-47,-4.84278e-47) (-5.1115e-48,-1.60718e-47) (-1.53538e-48,1.44548e-48) (1.35576e-48,2.98503e-48) (1.19873e-48,1.38946e-48) (5.9739e-49,4.69802e-49) (2.59055e-49,1.11572e-49) (9.37335e-50,-4.58545e-52) (2.30006e-50,-1.44951e-50) (2.28273e-51,-6.50885e-51) (-6.33027e-52,-1.41759e-51) (-2.97808e-52,-1.00867e-52) (-4.93713e-53,3.04048e-53) (-9.30423e-55,9.79009e-54) (1.18018e-54,9.99909e-55) (2.17408e-55,-6.55424e-56) (7.83544e-57,-3.02654e-56) (-2.9013e-57,-2.83059e-57) (-4.7072e-58,1.5262e-58) 
  (-3.34643e-62,7.88586e-63) (1.73428e-61,3.24173e-61) (2.68234e-60,-2.64381e-60) (-3.27654e-59,-1.71383e-59) (-5.09748e-59,3.42963e-58) (3.02709e-57,-6.46234e-58) (-1.4627e-56,-2.17702e-56) (-1.14284e-55,1.7657e-55) (1.57467e-54,2.3132e-55) (-3.42575e-54,-1.07979e-53) (-5.34157e-53,5.34568e-53) (4.5221e-52,1.29866e-52) (-6.83332e-52,-2.63249e-51) (-9.92619e-51,1.05783e-50) (6.99606e-50,1.12902e-50) (-1.40798e-49,-2.81175e-49) (-5.48306e-49,1.1291e-48) (4.3382e-48,-1.01716e-48) (-1.11917e-47,-8.26817e-48) (3.11873e-48,3.79148e-47) (6.25221e-47,-6.67645e-47) (-1.92514e-46,6.93963e-48) (2.72531e-46,1.98597e-46) (-1.98836e-46,-3.83447e-46) (1.68679e-46,2.8496e-46) (-4.37983e-46,2.97964e-47) (6.60086e-46,-3.07738e-46) (-2.44606e-46,5.48871e-46) (-5.6576e-46,-5.28528e-46) (8.53972e-46,-2.00679e-46) (-1.11446e-46,9.33243e-46) (-9.22527e-46,-4.08258e-46) (6.99689e-46,-7.46622e-46) (6.16801e-46,7.00573e-46) (-8.11648e-46,4.37493e-46) (-3.6681e-46,-6.82584e-46) (5.45927e-46,-3.53649e-46) (3.24953e-46,5.00572e-46) (-1.30223e-46,4.20474e-46) (-2.21324e-46,-1.24377e-46) (-1.47768e-46,-2.59117e-46) (-4.2281e-47,-7.7716e-47) (3.21426e-47,2.56187e-47) (3.63984e-47,1.09669e-47) (1.02153e-47,-1.00187e-47) (-3.10346e-48,-7.84511e-48) (-2.61624e-48,-1.67572e-48) (-1.64733e-49,2.4674e-49) (4.8597e-49,1.79045e-49) (3.18183e-49,1.19724e-50) (1.33911e-49,-2.4461e-50) (4.57137e-50,-2.19625e-50) (1.11602e-50,-1.26653e-50) (8.92099e-52,-4.84602e-51) (-5.73557e-52,-1.12332e-51) (-2.68544e-52,-1.00024e-52) (-5.26262e-53,2.57126e-53) (-2.68998e-54,1.05578e-53) (1.14808e-54,1.46696e-54) (2.94869e-55,-1.36963e-56) (2.23339e-56,-3.7488e-56) (-2.78961e-57,-5.36592e-57) (-7.88172e-58,-3.76987e-59) (-4.97422e-59,8.3176e-59) 
  (-5.62554e-63,5.11502e-63) (6.88232e-62,4.25951e-62) (2.03385e-61,-7.98157e-61) (-7.99578e-60,6.20454e-61) (3.0821e-59,6.78187e-59) (4.59638e-58,-4.712e-58) (-5.1256e-57,-2.04411e-57) (1.60001e-57,4.37356e-56) (2.9108e-55,-1.49951e-55) (-1.85854e-54,-1.36092e-54) (-2.17778e-54,1.50255e-53) (8.7004e-53,-3.38037e-53) (-4.21316e-52,-3.25537e-52) (-2.41813e-52,2.78938e-51) (1.17286e-50,-6.63016e-51) (-5.35799e-50,-2.42928e-50) (5.34482e-50,2.24559e-49) (4.88638e-49,-6.39745e-49) (-2.46924e-48,1.27242e-49) (4.63977e-48,4.79966e-48) (9.85577e-49,-1.58848e-47) (-2.43622e-47,2.23759e-47) (5.57884e-47,-5.81298e-48) (-6.39662e-47,-2.10903e-47) (4.69708e-47,4.80748e-48) (-4.21629e-47,6.48921e-47) (3.00145e-47,-1.11063e-46) (5.11471e-47,7.51163e-47) (-1.27147e-46,2.73365e-47) (5.08228e-47,-1.31809e-46) (1.17674e-46,1.01066e-46) (-1.43596e-46,8.79474e-47) (-3.48754e-47,-1.62434e-46) (1.56513e-46,-1.94684e-47) (-1.79971e-47,1.48524e-46) (-1.26906e-46,-1.38982e-47) (2.10993e-48,-1.08463e-46) (9.21664e-47,4.95305e-48) (4.51249e-47,6.30432e-47) (-3.05436e-47,1.74015e-47) (-4.70008e-47,-1.07574e-47) (-1.79252e-47,-4.21169e-48) (4.4792e-48,-3.84621e-49) (5.4527e-48,-2.5914e-48) (3.72809e-49,-2.39231e-48) (-1.20654e-48,-6.7503e-49) (-5.54818e-49,7.31315e-50) (-2.26395e-50,5.21156e-50) (7.16909e-50,-3.39946e-50) (3.84985e-50,-3.83142e-50) (1.25454e-50,-2.05907e-50) (2.42501e-51,-8.72927e-51) (-3.67012e-52,-3.00127e-51) (-5.34785e-52,-7.08695e-52) (-2.1982e-52,-6.47873e-53) (-4.7526e-53,2.24054e-53) (-3.53709e-54,1.02425e-53) (1.01459e-54,1.76173e-54) (3.46694e-55,5.07626e-56) (3.90468e-56,-4.0056e-56) (-1.70092e-57,-8.15145e-57) (-1.08872e-57,-4.05323e-58) (-1.18641e-58,9.58716e-59) (3.40167e-60,1.85392e-59) 
  (-5.08839e-64,1.59403e-63) (1.76882e-62,2.40194e-64) (-5.3913e-62,-1.70206e-61) (-1.37322e-60,1.03955e-60) (1.34138e-59,8.42251e-60) (2.44525e-59,-1.36323e-58) (-1.11908e-57,2.58553e-58) (5.47666e-57,7.15339e-57) (3.00935e-56,-5.94642e-56) (-4.6344e-55,1.80076e-57) (1.44947e-54,2.64713e-54) (9.52432e-54,-1.56518e-53) (-1.03125e-52,4.0709e-55) (2.94326e-52,4.46342e-52) (9.39983e-52,-2.35334e-51) (-1.05329e-50,2.76064e-51) (3.34107e-50,2.54553e-50) (-5.08827e-51,-1.43897e-49) (-3.22182e-49,2.93086e-49) (1.1554e-48,1.34748e-49) (-1.623e-48,-2.22002e-48) (-6.50647e-49,5.58544e-48) (6.11333e-48,-6.86117e-48) (-9.17108e-48,4.59856e-48) (4.24e-48,-5.25121e-48) (4.29729e-48,1.27505e-47) (-1.0171e-47,-1.44658e-47) (1.40417e-47,-1.025e-48) (-8.57233e-48,1.98276e-47) (-1.29747e-47,-1.8535e-47) (2.46279e-47,-6.748e-48) (-1.67575e-48,2.78131e-47) (-2.47836e-47,-1.01716e-47) (1.23102e-47,-2.34215e-47) (1.79017e-47,1.60527e-47) (-1.3656e-47,1.5795e-47) (-1.46166e-47,-1.05166e-47) (8.67538e-48,-1.10831e-47) (1.32742e-47,6.28122e-49) (3.05875e-49,5.00115e-48) (-6.19945e-48,4.29393e-48) (-2.95431e-48,1.98835e-48) (2.39815e-49,-2.43385e-49) (3.52057e-49,-8.53646e-49) (-1.95068e-49,-3.55333e-49) (-2.20852e-49,3.80832e-50) (-6.614e-50,7.33301e-50) (-2.84516e-52,1.28277e-50) (3.73766e-51,-1.1112e-50) (-3.05234e-52,-9.10146e-51) (-1.21699e-51,-4.04123e-51) (-8.78255e-52,-1.34537e-51) (-4.42859e-52,-3.06368e-52) (-1.58335e-52,-1.49522e-53) (-3.5745e-53,2.08463e-53) (-3.10556e-54,9.053e-54) (8.73286e-55,1.78953e-54) (3.62742e-55,1.01822e-55) (5.3329e-56,-3.7952e-56) (1.94432e-58,-1.05257e-56) (-1.28459e-57,-9.16588e-58) (-2.05742e-58,8.23719e-59) (-4.70957e-60,2.8902e-59) (2.86094e-60,2.25143e-60) 
  (8.33778e-65,3.55765e-64) (3.28554e-63,-1.97056e-63) (-2.93912e-62,-2.45809e-62) (-1.22991e-61,3.4473e-61) (3.33006e-60,-1.0337e-61) (-1.18856e-59,-2.62632e-59) (-1.57932e-58,1.76045e-58) (1.7554e-57,5.34065e-58) (-2.1733e-57,-1.32446e-56) (-7.37924e-56,5.53779e-56) (5.41701e-55,2.42837e-55) (-3.90426e-55,-3.53727e-54) (-1.55126e-53,1.22472e-53) (9.60069e-53,3.14251e-53) (-1.38367e-52,-4.50863e-52) (-1.17744e-51,1.60944e-51) (7.5599e-51,-2.64899e-52) (-1.6862e-50,-1.91415e-50) (-1.11457e-50,7.52865e-50) (1.69448e-49,-1.08761e-49) (-4.57837e-49,-1.13472e-49) (5.34714e-49,7.79787e-49) (-2.48857e-50,-1.48124e-48) (-4.66626e-49,1.44972e-48) (-3.64891e-49,-9.32004e-49) (2.14234e-48,8.15688e-49) (-2.6351e-48,-1.83458e-49) (9.67607e-49,-2.04654e-48) (1.80014e-48,3.04131e-48) (-3.61499e-48,9.18603e-50) (1.35907e-48,-3.96166e-48) (3.56836e-48,2.84867e-48) (-3.58491e-48,2.37688e-48) (-1.99357e-48,-3.91767e-48) (3.73025e-48,-8.90821e-49) (8.47848e-49,3.283e-48) (-2.80062e-48,9.69222e-49) (-6.68628e-49,-2.02499e-48) (1.47307e-48,-1.65304e-48) (7.37848e-49,2.61397e-49) (-1.45624e-49,1.13055e-48) (-1.06766e-49,6.43393e-49) (9.07722e-51,1.00856e-50) (-4.51739e-50,-1.2753e-49) (-6.1519e-50,-2.58562e-50) (-2.37449e-50,2.7006e-50) (-4.16862e-52,1.70949e-50) (1.43515e-51,2.44831e-51) (-7.84061e-52,-1.45915e-51) (-1.13417e-51,-9.8208e-52) (-6.59981e-52,-3.11301e-52) (-2.79644e-52,-4.10147e-53) (-9.26329e-53,2.25006e-53) (-2.09651e-53,1.90429e-53) (-1.66392e-54,7.23705e-54) (7.87451e-55,1.54288e-54) (3.44164e-55,1.1698e-55) (6.0745e-56,-3.34668e-56) (2.24435e-57,-1.19354e-56) (-1.32415e-57,-1.45565e-57) (-2.94604e-58,3.78916e-59) (-1.82836e-59,3.78002e-59) (3.01425e-60,4.69986e-60) (6.97222e-61,-4.04882e-62) 
  (5.57311e-65,5.60537e-65) (3.68628e-64,-7.33935e-64) (-8.07781e-63,-9.6856e-64) (1.87136e-62,7.46354e-62) (5.60237e-61,-4.08325e-61) (-5.0996e-60,-3.0378e-60) (-5.45131e-60,4.78722e-59) (3.49645e-58,-1.20288e-58) (-1.91481e-57,-1.86762e-57) (-5.08387e-57,1.74509e-56) (1.12514e-55,-2.63622e-56) (-4.75848e-55,-4.91449e-55) (-8.75878e-55,3.64481e-54) (1.76975e-53,-6.60042e-54) (-7.19796e-53,-4.86115e-53) (1.8722e-53,3.60957e-52) (1.01324e-51,-8.90257e-52) (-4.41951e-51,-7.25607e-52) (6.76369e-51,1.13352e-50) (1.06371e-50,-3.29529e-50) (-7.2009e-50,3.54557e-50) (1.52323e-49,3.84954e-50) (-1.62875e-49,-1.69041e-49) (1.04922e-49,1.93016e-49) (-1.58152e-49,-1.86863e-50) (3.33802e-49,-1.84315e-49) (-2.56236e-49,2.84967e-49) (-2.13327e-49,-3.11001e-49) (5.65601e-49,5.55117e-50) (-3.04946e-49,4.91872e-49) (-4.06859e-49,-5.49141e-49) (7.11512e-49,-2.05501e-49) (-4.56734e-51,6.89208e-49) (-7.13412e-49,-1.09511e-49) (2.17734e-49,-5.68013e-49) (5.13009e-49,1.89421e-49) (-1.37356e-49,4.62181e-49) (-3.14683e-49,-7.89755e-50) (-5.56626e-50,-3.5417e-49) (9.46801e-50,-9.78763e-50) (1.0943e-49,1.24962e-49) (6.86772e-50,9.13537e-50) (1.07318e-50,6.60656e-51) (-1.64276e-50,-9.18074e-51) (-1.03166e-50,3.01278e-51) (-2.45847e-52,5.70637e-51) (1.84746e-51,2.24769e-51) (5.45198e-52,2.34073e-52) (-2.14688e-52,-5.10208e-53) (-2.41211e-52,2.76407e-53) (-1.14954e-52,4.80212e-53) (-3.77291e-53,3.17168e-53) (-7.88594e-54,1.47956e-53) (-4.28067e-57,5.01385e-54) (7.40049e-55,1.0985e-54) (2.98162e-55,9.02981e-56) (5.8955e-56,-2.95083e-56) (3.59564e-57,-1.21621e-56) (-1.23236e-57,-1.86853e-57) (-3.64376e-58,-2.68821e-59) (-3.54727e-59,4.2728e-59) (2.26871e-60,7.56971e-60) (1.02008e-60,2.78525e-61) (9.41475e-62,-9.40533e-62) 
  (1.64954e-65,3.77281e-66) (-1.89886e-65,-1.73148e-64) (-1.5265e-63,7.67932e-64) (1.19273e-62,1.06661e-62) (4.70502e-62,-1.3472e-61) (-1.20569e-60,9.26803e-62) (4.73456e-60,8.48042e-60) (4.21562e-59,-6.05003e-59) (-5.22833e-58,-7.04656e-59) (1.25963e-57,3.31281e-57) (1.41065e-56,-1.72262e-56) (-1.28877e-55,-1.81197e-56) (2.95175e-55,6.38746e-55) (1.79387e-54,-2.99986e-54) (-1.57736e-53,1.36059e-54) (4.3514e-53,4.80838e-53) (3.90184e-53,-2.34972e-52) (-6.75771e-52,3.88897e-52) (2.13704e-51,7.75608e-52) (-2.18159e-51,-5.49955e-51) (-5.37822e-51,1.24269e-50) (2.28686e-50,-1.18964e-50) (-3.64726e-50,-1.77082e-51) (2.97852e-50,7.38927e-51) (-1.6052e-50,2.19219e-50) (1.26801e-50,-6.04784e-50) (1.10713e-50,5.29466e-50) (-6.40608e-50,2.80295e-51) (5.98255e-50,-6.69336e-50) (3.93428e-50,8.42234e-50) (-1.10734e-49,3.35505e-51) (3.91688e-50,-1.12265e-49) (9.12912e-50,6.20743e-50) (-8.22982e-50,8.31485e-50) (-5.49507e-50,-7.88911e-50) (7.18533e-50,-5.01398e-50) (4.70832e-50,6.14076e-50) (-3.57303e-50,3.51486e-50) (-4.86034e-50,-2.86531e-50) (-7.21367e-51,-2.39237e-50) (2.3245e-50,-3.02522e-52) (1.91409e-50,2.29916e-51) (3.63099e-51,-6.83723e-52) (-2.40376e-51,4.56063e-52) (-9.48049e-52,1.39408e-51) (5.33003e-52,7.21908e-52) (4.80049e-52,8.14051e-53) (1.13601e-52,-3.16529e-53) (-2.12497e-53,1.68022e-53) (-2.25e-53,3.13446e-53) (-6.97591e-54,1.98051e-53) (-2.4525e-55,8.5131e-54) (1.01064e-54,2.74861e-54) (6.52432e-55,5.93782e-55) (2.31919e-55,3.67948e-56) (4.85131e-56,-2.73289e-56) (3.65332e-57,-1.13054e-56) (-1.09419e-57,-2.02778e-57) (-4.0028e-58,-8.79799e-59) (-5.20699e-59,4.2782e-59) (6.12677e-61,1.0296e-59) (1.27043e-60,7.54051e-61) (1.77398e-61,-9.00273e-62) (1.4315e-63,-2.51489e-62) 
  (3.3684e-66,-1.22204e-66) (-2.33182e-65,-2.81316e-65) (-1.73967e-64,3.09452e-64) (3.2646e-63,4.19927e-64) (-7.87491e-63,-2.79735e-62) (-1.87144e-61,1.5619e-61) (1.75731e-60,8.16128e-61) (-3.79929e-61,-1.45496e-59) (-8.99686e-59,5.01333e-59) (5.80461e-58,3.61981e-58) (1.23193e-58,-4.24459e-57) (-2.1215e-56,1.22719e-56) (1.16719e-55,5.89025e-56) (-8.76157e-56,-6.34212e-55) (-2.05716e-54,1.98213e-54) (1.13889e-53,1.73859e-54) (-2.07139e-53,-3.61665e-53) (-4.80129e-53,1.25815e-52) (3.6716e-52,-1.28526e-52) (-8.8091e-52,-4.81942e-52) (6.70878e-52,2.16132e-51) (1.46607e-51,-3.90661e-51) (-4.21365e-51,3.64054e-51) (3.37397e-51,-2.39286e-51) (1.7365e-51,4.47732e-51) (-5.88414e-51,-7.76324e-51) (6.9506e-51,2.77998e-51) (-5.68356e-51,9.33372e-51) (-2.97948e-51,-1.362e-50) (1.48373e-50,2.15953e-51) (-9.78068e-51,1.48917e-50) (-1.09619e-50,-1.54014e-50) (1.6411e-50,-6.5937e-51) (2.97558e-51,1.84696e-50) (-1.51633e-50,2.23527e-52) (3.60728e-54,-1.39469e-50) (1.22324e-50,-2.86216e-52) (1.83824e-51,7.70118e-51) (-8.09968e-51,2.98096e-51) (-4.38417e-51,-1.32105e-51) (1.91606e-51,-2.44937e-51) (2.42991e-51,-1.99011e-51) (4.8792e-52,-6.86018e-52) (-1.95335e-52,2.13351e-52) (2.44165e-53,2.55255e-52) (1.34783e-52,3.49154e-53) (6.83968e-53,-4.1873e-53) (1.26639e-53,-1.85898e-53) (4.44196e-55,2.95877e-54) (1.31814e-54,5.87449e-54) (1.67155e-54,3.06785e-54) (1.05861e-54,1.00174e-54) (4.72109e-55,1.87024e-55) (1.53543e-55,-1.4694e-56) (3.25653e-56,-2.5525e-56) (2.43339e-57,-9.58666e-57) (-9.90015e-58,-1.88332e-57) (-3.98431e-58,-1.19443e-58) (-6.32678e-59,3.94431e-59) (-1.46842e-60,1.22619e-59) (1.38377e-60,1.30659e-60) (2.68331e-61,-5.73444e-62) (1.31962e-62,-3.47601e-62) (-2.9575e-63,-3.70005e-63) 
  (4.4927e-67,-6.01112e-67) (-7.26753e-66,-2.15875e-66) (6.3101e-66,7.26826e-65) (5.94419e-64,-3.08879e-64) (-4.54938e-63,-3.6875e-63) (-1.21368e-62,4.70897e-62) (3.75268e-61,-7.44718e-62) (-1.75306e-60,-2.23911e-60) (-8.0613e-60,1.81997e-59) (1.30125e-58,-1.24019e-59) (-4.72702e-58,-6.47574e-58) (-1.6957e-57,4.24279e-57) (2.3545e-56,-4.89043e-57) (-8.44535e-56,-7.96608e-56) (-6.24645e-56,5.06511e-55) (1.74699e-54,-1.02842e-54) (-6.74863e-54,-2.59267e-54) (7.23629e-54,2.19253e-53) (3.44811e-53,-5.64476e-53) (-1.65999e-52,3.28228e-53) (3.18073e-52,1.97504e-52) (-2.45579e-52,-6.18851e-52) (-7.56325e-53,8.27579e-52) (2.45869e-53,-5.36687e-52) (8.22283e-52,2.12507e-52) (-1.48815e-51,-1.00268e-52) (8.16368e-52,-6.40404e-52) (7.25034e-52,1.6931e-51) (-1.96526e-51,-8.32242e-52) (1.62194e-51,-1.80217e-51) (1.04086e-51,2.64252e-51) (-2.97891e-51,9.99173e-54) (5.99409e-52,-2.76819e-51) (2.6286e-51,1.34145e-51) (-1.30591e-51,2.0013e-51) (-1.80538e-51,-1.26658e-51) (1.08754e-51,-1.56508e-51) (1.21331e-51,3.99716e-52) (-4.09398e-52,1.21667e-51) (-6.55746e-52,4.87622e-52) (-1.10425e-52,-3.80607e-52) (3.87408e-53,-4.93535e-52) (-2.65139e-53,-1.67977e-52) (-7.52792e-54,2.89923e-53) (2.66035e-53,2.65941e-53) (1.93331e-53,-8.89624e-54) (3.86026e-54,-1.24189e-53) (-4.87625e-55,-4.11893e-54) (3.41237e-55,-2.22372e-57) (8.12362e-55,4.37341e-55) (5.58477e-55,1.31961e-55) (2.46084e-55,-2.05812e-56) (7.81626e-56,-3.90601e-56) (1.60281e-56,-2.14705e-56) (5.97482e-58,-7.22135e-57) (-9.31293e-58,-1.47703e-57) (-3.63065e-58,-1.0757e-58) (-6.56297e-59,3.54982e-59) (-3.16564e-60,1.30996e-59) (1.35541e-60,1.79413e-60) (3.48912e-61,-7.90871e-65) (2.90823e-62,-4.14493e-62) (-2.54611e-63,-6.41752e-63) (-8.7322e-64,-1.43745e-64) 
  (8.38597e-69,-1.55228e-67) (-1.48314e-66,4.70726e-67) (9.45102e-66,1.14331e-65) (6.22456e-65,-1.19686e-64) (-1.16571e-63,-7.1868e-65) (3.5145e-63,8.93624e-63) (5.04648e-62,-5.51904e-62) (-5.30845e-61,-1.44201e-61) (8.73314e-61,3.70736e-60) (1.80915e-59,-1.686e-59) (-1.44102e-58,-4.11994e-59) (2.39342e-58,8.0867e-58) (2.79585e-57,-3.37056e-57) (-2.07806e-56,-1.62482e-57) (4.78691e-56,7.65563e-56) (1.23061e-55,-3.31317e-55) (-1.18212e-54,3.86786e-55) (3.31211e-54,2.11843e-54) (-1.54729e-54,-1.10705e-53) (-1.77053e-53,2.20759e-53) (6.04564e-53,-9.95564e-54) (-9.41365e-53,-4.56757e-53) (7.64061e-53,9.39526e-53) (-5.48598e-53,-4.0016e-53) (1.16981e-52,-8.96586e-53) (-1.55549e-52,1.57566e-52) (-3.01106e-53,-1.46832e-52) (2.96158e-52,7.11471e-53) (-2.72637e-52,1.74089e-52) (-9.32158e-53,-3.80594e-52) (4.35643e-52,1.07063e-52) (-2.66782e-52,3.81798e-52) (-3.10752e-52,-3.29233e-52) (4.09938e-52,-2.07452e-52) (1.45973e-52,3.46814e-52) (-3.25869e-52,1.17202e-52) (-9.64497e-53,-2.76265e-52) (1.62334e-52,-1.31187e-52) (1.02348e-52,1.55063e-52) (-4.68407e-54,1.40933e-52) (-4.71584e-53,-1.18958e-53) (-5.03391e-53,-5.62807e-53) (-2.56373e-53,-1.89168e-53) (-6.79774e-55,3.08479e-54) (5.25595e-54,5.56514e-55) (1.39094e-54,-2.8745e-54) (-8.50424e-55,-1.8943e-54) (-5.55402e-55,-4.93949e-55) (-7.96127e-58,-6.88939e-56) (1.29087e-55,-5.15676e-56) (7.62067e-56,-5.34289e-56) (2.49337e-56,-3.30733e-56) (3.93831e-57,-1.43862e-56) (-8.87158e-58,-4.53695e-57) (-8.52206e-58,-9.29492e-58) (-3.0055e-58,-5.94635e-59) (-5.83601e-59,3.28639e-59) (-3.74771e-60,1.27627e-59) (1.24758e-60,2.07452e-60) (4.01933e-61,6.29221e-62) (4.60954e-62,-4.37642e-62) (-1.28492e-63,-9.19496e-63) (-1.14683e-63,-5.54549e-64) (-1.38105e-64,8.89709e-65) 
  (-1.63751e-68,-2.73237e-68) (-1.9424e-67,2.4923e-67) (2.87556e-66,7.99063e-67) (-3.66518e-66,-2.66378e-65) (-1.95116e-64,1.22843e-64) (1.58486e-63,1.00604e-63) (1.49246e-63,-1.43962e-62) (-9.78843e-62,3.898e-62) (5.57271e-61,4.58552e-61) (7.52412e-61,-4.57129e-60) (-2.57087e-59,1.04264e-59) (1.26029e-58,8.87338e-59) (1.40331e-59,-7.8954e-58) (-3.05713e-57,2.09491e-57) (1.4967e-56,5.135e-57) (-1.96091e-56,-5.78443e-56) (-1.15016e-55,1.78503e-55) (6.60915e-55,-7.56907e-56) (-1.38309e-54,-1.26927e-54) (1.30479e-55,4.69205e-54) (6.26313e-54,-7.68103e-54) (-1.54867e-53,4.68656e-54) (1.7084e-53,1.81735e-54) (-7.788e-54,3.96487e-54) (9.46659e-55,-2.4877e-53) (2.85526e-54,3.16627e-53) (-2.28079e-53,-5.4725e-54) (3.82513e-53,-3.09913e-53) (-8.57241e-55,4.88604e-53) (-5.88272e-53,-2.26947e-53) (5.31099e-53,-4.59361e-53) (2.47986e-53,6.79661e-53) (-7.12844e-53,1.06688e-53) (1.11827e-53,-6.97659e-53) (5.80016e-53,1.17114e-53) (-1.44404e-53,5.20074e-53) (-4.25599e-53,-1.25103e-53) (-2.81726e-54,-3.40304e-53) (2.61868e-53,1.49555e-54) (1.75681e-53,1.56256e-53) (-3.60673e-54,4.98539e-54) (-1.11285e-53,-3.28381e-55) (-5.5922e-54,8.1723e-55) (-2.04072e-55,6.38352e-55) (6.00725e-55,-3.67928e-55) (-1.12382e-55,-4.5448e-55) (-2.97755e-55,-1.33503e-55) (-1.29921e-55,8.9799e-58) (-1.59633e-56,-6.79815e-57) (5.96622e-57,-1.97732e-56) (1.64857e-57,-1.48184e-56) (-1.34067e-57,-6.7446e-57) (-1.36852e-57,-2.12209e-57) (-6.7811e-58,-4.09331e-58) (-2.18065e-58,-6.86966e-61) (-4.35072e-59,3.10086e-59) (-2.97027e-60,1.13934e-59) (1.14213e-60,2.06145e-60) (4.18859e-61,1.06299e-61) (5.97237e-62,-4.22343e-62) (5.73174e-64,-1.14924e-62) (-1.3164e-63,-1.0625e-63) (-2.23506e-64,6.77852e-65) (-7.81728e-66,2.9279e-65) 
  (-5.86583e-69,-2.70254e-69) (-3.54345e-69,6.33991e-68) (5.59868e-67,-1.99454e-67) (-3.64315e-66,-3.85664e-66) (-1.67945e-65,4.1818e-65) (3.62525e-64,-2.47318e-65) (-1.41908e-63,-2.38331e-63) (-1.0359e-62,1.70901e-62) (1.35334e-61,4.76267e-63) (-4.09401e-61,-7.55724e-61) (-2.52663e-60,4.41333e-60) (2.78503e-59,-1.60385e-60) (-8.62211e-59,-1.11588e-58) (-1.87169e-58,6.25245e-58) (2.58044e-57,-9.44125e-58) (-8.85583e-57,-5.57961e-57) (3.92156e-57,3.57821e-56) (7.81285e-56,-8.00769e-56) (-3.12824e-55,-1.57388e-56) (5.18029e-55,5.71948e-55) (-6.95609e-56,-1.58192e-54) (-1.23733e-54,2.12564e-54) (1.82783e-54,-1.49815e-54) (1.26224e-55,1.25628e-54) (-2.9914e-54,-2.77648e-54) (3.64889e-54,2.46469e-54) (-2.5705e-54,3.01007e-54) (-1.53172e-55,-7.76313e-54) (6.17007e-54,4.11709e-54) (-8.39715e-54,5.55105e-54) (-1.05508e-54,-1.08476e-53) (1.08045e-53,2.86531e-54) (-5.13115e-54,1.01856e-53) (-7.62861e-54,-7.57263e-54) (6.67018e-54,-6.45452e-54) (5.25862e-54,6.47983e-54) (-5.21361e-54,4.14112e-54) (-4.76009e-54,-2.83511e-54) (2.24325e-54,-2.85883e-54) (3.75626e-54,-5.19331e-55) (5.7882e-55,7.28633e-55) (-1.11628e-54,1.12209e-54) (-5.75528e-55,7.678e-55) (1.7931e-56,1.68151e-55) (3.59121e-56,-8.03751e-56) (-5.37708e-56,-3.93388e-56) (-4.80208e-56,1.54247e-56) (-1.62933e-56,1.50945e-56) (-3.40226e-57,2.03756e-57) (-1.80734e-57,-2.45179e-57) (-1.59936e-57,-1.73652e-57) (-9.74639e-58,-5.7208e-58) (-4.18606e-58,-6.66356e-59) (-1.29045e-58,3.87612e-59) (-2.54677e-59,2.7478e-59) (-1.25122e-60,9.17412e-60) (1.07489e-60,1.75408e-60) (3.99833e-61,1.11169e-61) (6.59757e-62,-3.90566e-62) (2.36877e-63,-1.28547e-62) (-1.35556e-63,-1.56469e-63) (-3.05449e-64,2.32638e-65) (-2.14881e-65,3.67326e-65) (2.55943e-66,4.93065e-66) 
  (-1.27673e-69,2.21902e-70) (6.6512e-69,1.0737e-68) (6.72578e-68,-9.5941e-68) (-1.01774e-66,-1.95855e-67) (2.14392e-66,8.45421e-66) (5.30595e-65,-4.51289e-65) (-4.86815e-64,-2.00495e-64) (3.91432e-64,3.73387e-63) (2.04773e-62,-1.46307e-62) (-1.44664e-61,-6.33556e-62) (1.35406e-61,9.13271e-61) (3.72732e-60,-3.3336e-60) (-2.42484e-59,-5.84685e-60) (4.31291e-59,1.05386e-58) (2.42851e-58,-4.05839e-58) (-1.76713e-57,2.10777e-58) (4.3073e-57,4.26504e-57) (1.64671e-57,-1.86317e-56) (-4.14651e-56,3.12185e-56) (1.24719e-55,1.53114e-56) (-1.74942e-55,-1.7818e-55) (8.25209e-56,3.57669e-55) (2.40542e-56,-3.12491e-55) (2.05009e-55,6.22793e-56) (-6.45552e-55,6.57319e-56) (5.56604e-55,-1.86678e-55) (2.232e-55,6.53728e-55) (-9.5641e-55,-7.15916e-55) (1.04013e-54,-4.6552e-55) (-6.8091e-56,1.58828e-54) (-1.45888e-54,-8.31115e-55) (1.31096e-54,-1.11279e-54) (8.29917e-55,1.58593e-54) (-1.59676e-54,2.77717e-55) (-2.31599e-55,-1.43138e-54) (1.27679e-54,-7.90993e-56) (6.6521e-56,9.90822e-55) (-8.17299e-55,3.41104e-55) (-1.66585e-55,-4.72081e-55) (3.2259e-55,-4.9668e-55) (1.62404e-55,-5.19059e-56) (9.62251e-57,2.15749e-55) (2.20033e-56,1.55354e-55) (2.48869e-56,2.78147e-56) (-6.23514e-58,-1.03076e-56) (-9.0946e-57,6.12234e-58) (-3.81538e-57,6.64089e-57) (-2.87264e-58,3.70906e-57) (-1.38097e-58,8.15655e-58) (-4.51012e-58,1.28874e-59) (-3.69591e-58,1.36106e-59) (-1.74815e-58,5.70377e-59) (-5.47273e-59,4.45158e-59) (-9.76796e-60,2.05491e-59) (5.10315e-61,6.37386e-60) (1.00499e-60,1.23806e-60) (3.4907e-61,7.60244e-62) (6.28719e-62,-3.63746e-62) (3.35943e-63,-1.30961e-62) (-1.29744e-63,-1.92514e-63) (-3.68659e-64,-3.36203e-65) (-3.70736e-65,4.08056e-65) (1.68073e-66,7.52096e-66) (9.50707e-67,3.47229e-67) 
  (-1.82961e-70,1.81027e-70) (2.28899e-69,9.72956e-70) (-2.11249e-70,-2.28706e-68) (-1.81673e-67,8.48303e-68) (1.29021e-66,1.06316e-66) (2.97086e-66,-1.28875e-65) (-9.57851e-65,2.49582e-65) (4.79323e-64,5.08264e-64) (1.33737e-63,-4.43577e-63) (-2.78471e-62,7.12496e-63) (1.20906e-61,1.13784e-61) (1.48429e-61,-8.75416e-61) (-3.95415e-60,1.86254e-60) (1.72481e-59,9.49249e-60) (-1.13414e-59,-7.99216e-59) (-2.09505e-58,2.15239e-58) (1.00946e-57,1.00548e-58) (-1.75194e-57,-2.56815e-57) (-1.91333e-57,8.32045e-57) (1.67721e-56,-1.1352e-56) (-3.87739e-56,-2.26018e-57) (4.47446e-56,2.97006e-56) (-2.71867e-56,-2.89783e-56) (2.8207e-56,-2.72357e-56) (-5.85458e-56,8.10756e-56) (2.06604e-56,-7.26468e-56) (1.1592e-55,3.14075e-56) (-1.7291e-55,4.79717e-56) (2.49375e-56,-1.76068e-55) (1.93372e-55,1.55079e-55) (-2.32584e-55,1.09442e-55) (-2.53894e-56,-2.62351e-55) (2.75241e-55,4.03968e-56) (-1.02991e-55,2.19856e-55) (-2.02337e-55,-9.88597e-56) (1.03051e-55,-1.64783e-55) (1.27695e-55,7.44709e-56) (-3.52153e-56,1.34376e-55) (-6.90173e-56,-1.26861e-56) (-2.4683e-56,-8.617e-56) (6.69165e-57,-3.19536e-56) (2.17936e-56,1.76885e-56) (1.98194e-56,1.48992e-56) (7.35076e-57,1.07175e-57) (-3.81929e-58,-1.20293e-57) (-8.51828e-58,8.17065e-58) (2.54445e-58,1.11192e-57) (3.81931e-58,4.77277e-58) (9.94092e-59,1.27542e-58) (-3.53277e-59,5.84686e-59) (-3.52362e-59,4.53238e-59) (-1.17046e-59,2.72216e-59) (-5.37713e-61,1.16277e-59) (1.45707e-60,3.52387e-60) (8.54509e-61,6.6694e-61) (2.7222e-61,1.91493e-62) (5.11047e-62,-3.45006e-62) (3.11012e-63,-1.22477e-62) (-1.21059e-63,-2.03729e-63) (-4.01637e-64,-8.15722e-65) (-5.12786e-65,4.12274e-65) (2.16058e-67,9.86001e-66) (1.14511e-66,7.82807e-67) (1.69257e-67,-7.03145e-68) 
  (-9.00897e-72,4.98064e-71) (4.73758e-70,-1.03865e-70) (-2.61601e-69,-3.56467e-69) (-1.85541e-68,3.36417e-68) (3.1698e-67,1.68954e-68) (-1.00384e-66,-2.27598e-66) (-1.14193e-65,1.4473e-65) (1.27126e-64,2.06389e-65) (-3.02856e-64,-7.88767e-64) (-3.15903e-63,4.10853e-63) (2.94692e-62,2.52081e-63) (-7.56967e-62,-1.36623e-61) (-3.32505e-61,6.82197e-61) (3.32218e-60,-5.90224e-61) (-9.99736e-60,-9.31994e-60) (-4.64181e-60,5.01344e-59) (1.4096e-58,-9.2844e-59) (-4.93204e-58,-1.43322e-58) (6.40311e-58,1.23739e-57) (8.12023e-58,-3.12512e-57) (-4.62265e-57,3.753e-57) (7.5693e-57,-1.34881e-57) (-4.75195e-57,2.52457e-58) (-1.15057e-57,-7.03454e-57) (3.21792e-57,1.4577e-56) (-6.71194e-57,-6.81115e-57) (1.59987e-56,-1.26871e-56) (-9.68645e-57,2.45149e-56) (-2.12961e-56,-1.83812e-56) (3.68523e-56,-9.73612e-57) (-6.69855e-57,3.85778e-56) (-3.51134e-56,-1.97124e-56) (3.00162e-56,-3.04611e-56) (1.82803e-56,3.12793e-56) (-3.0542e-56,1.64996e-56) (-1.11604e-56,-2.70516e-56) (1.98128e-56,-9.68841e-57) (1.29854e-56,1.69289e-56) (-6.4032e-57,8.04504e-57) (-1.19223e-56,-5.54076e-57) (-4.10635e-57,-4.43189e-57) (3.36858e-57,-6.6312e-58) (3.75439e-57,-5.39376e-58) (1.14838e-57,-7.5783e-58) (-8.80235e-59,-1.93717e-58) (-1.66877e-59,1.39515e-58) (1.38218e-58,9.23635e-59) (9.7689e-59,1.35202e-59) (2.99958e-59,2.86233e-60) (4.93115e-60,9.55795e-60) (1.96315e-60,8.62853e-60) (2.04596e-60,4.26557e-60) (1.36196e-60,1.33083e-60) (5.97463e-61,2.12804e-61) (1.79983e-61,-3.02078e-62) (3.3962e-62,-3.16203e-62) (1.75947e-63,-1.04295e-62) (-1.14361e-63,-1.86195e-63) (-4.00533e-64,-1.003e-64) (-6.01927e-65,3.93606e-65) (-1.43072e-66,1.15364e-65) (1.23765e-66,1.24246e-66) (2.45246e-67,-3.80096e-68) (1.37844e-68,-2.99726e-68) 
  (4.165e-72,8.93397e-72) (6.27514e-71,-6.95496e-71) (-8.0612e-70,-2.59011e-70) (9.35708e-70,7.23236e-69) (4.97724e-68,-3.29845e-68) (-4.043e-67,-2.26732e-67) (-6.10809e-68,3.40132e-66) (2.07023e-65,-1.11685e-65) (-1.30694e-64,-7.88915e-65) (9.91174e-66,9.25726e-64) (4.35105e-63,-2.88433e-63) (-2.51759e-62,-1.03601e-62) (2.8957e-62,1.27348e-61) (3.76612e-61,-4.32436e-61) (-2.29098e-60,-1.64347e-61) (4.64413e-60,6.98288e-60) (8.40083e-60,-2.66328e-59) (-7.73441e-59,3.35796e-59) (2.0889e-58,8.47469e-59) (-2.31198e-58,-4.53342e-58) (-1.29982e-58,8.89541e-58) (6.30717e-58,-8.69732e-58) (-2.85684e-58,4.47922e-58) (-1.09499e-57,-6.03996e-58) (1.88337e-57,1.04753e-57) (-1.18141e-57,4.60583e-58) (-2.47521e-59,-3.37214e-57) (2.03339e-57,3.211e-57) (-4.31971e-57,1.19813e-57) (2.13791e-57,-5.36927e-57) (4.21089e-57,4.19049e-57) (-5.52217e-57,2.66397e-57) (-1.01923e-57,-6.41755e-57) (5.38694e-57,3.75485e-58) (-6.93556e-58,5.25795e-57) (-4.25487e-57,-9.88066e-58) (4.29958e-58,-3.27967e-57) (3.20556e-57,3.08759e-59) (6.27664e-58,1.4645e-57) (-1.69908e-57,7.75373e-58) (-1.06252e-57,7.93056e-59) (1.63463e-58,-3.52513e-58) (3.34789e-58,-4.51115e-58) (5.79693e-59,-2.34434e-58) (-3.14753e-59,-3.25821e-59) (7.2733e-60,1.24143e-59) (2.32476e-59,-4.26652e-60) (1.26506e-59,-9.17958e-60) (4.10053e-60,-3.52769e-60) (1.76593e-60,1.36833e-61) (1.22307e-60,5.90938e-61) (7.22605e-61,1.96487e-61) (3.08103e-61,-2.1989e-62) (9.20978e-62,-4.97593e-62) (1.6583e-62,-2.56132e-62) (-3.36064e-67,-7.83952e-63) (-1.08294e-63,-1.44168e-63) (-3.66623e-64,-8.15032e-65) (-6.11205e-65,3.71249e-65) (-2.61708e-66,1.22698e-65) (1.23386e-66,1.62665e-66) (3.09908e-67,7.34498e-69) (2.71166e-68,-3.48277e-68) (-1.84014e-69,-5.6089e-69) 
  (1.65368e-72,9.38591e-73) (1.97154e-72,-1.78138e-71) (-1.52548e-70,5.0323e-71) (9.48706e-70,9.90457e-70) (3.76033e-69,-1.04741e-68) (-8.48046e-68,1.15515e-68) (3.68494e-67,5.01105e-67) (1.73054e-66,-3.88942e-66) (-2.71353e-65,3.25867e-66) (1.02789e-64,1.27611e-64) (2.81889e-64,-8.68368e-64) (-4.51379e-63,1.31947e-63) (1.74598e-62,1.38408e-62) (3.7375e-63,-9.66045e-62) (-3.14945e-61,2.18442e-61) (1.32464e-60,4.16523e-61) (-1.69991e-60,-4.26886e-60) (-6.16866e-60,1.22886e-59) (3.42278e-59,-1.1603e-59) (-7.38952e-59,-2.86035e-59) (7.56365e-59,1.10072e-58) (-2.10975e-59,-1.44492e-58) (2.96941e-59,4.77781e-59) (-1.96793e-58,7.53513e-59) (2.82258e-58,-1.02085e-58) (4.2829e-60,1.9239e-58) (-4.22657e-58,-3.36478e-58) (5.40959e-58,2.29928e-59) (-2.3603e-58,6.73649e-58) (-4.5682e-58,-7.33952e-58) (8.84398e-58,-1.57604e-58) (-1.5085e-58,9.17625e-58) (-8.65816e-58,-4.49708e-58) (4.97088e-58,-6.34079e-58) (5.80293e-58,5.5378e-58) (-4.84029e-58,4.29149e-58) (-3.75902e-58,-3.28242e-58) (2.93605e-58,-3.68469e-58) (2.55262e-58,3.17437e-59) (-6.77795e-59,2.47601e-58) (-1.05661e-58,1.45155e-58) (-2.49879e-59,-3.1968e-59) (-1.23769e-59,-7.9506e-59) (-1.99222e-59,-3.53647e-59) (-9.17434e-60,-2.41986e-60) (8.56568e-61,5.78094e-61) (1.84167e-60,-2.69682e-60) (4.11828e-61,-2.39914e-60) (5.48861e-62,-9.40201e-61) (1.8405e-61,-2.39484e-61) (1.8677e-61,-9.24426e-62) (9.72e-62,-6.62212e-62) (3.0156e-62,-3.9498e-62) (4.02027e-63,-1.66674e-62) (-1.28455e-63,-4.90021e-63) (-9.64155e-64,-8.95381e-64) (-3.03504e-64,-3.46574e-65) (-5.35217e-65,3.53891e-65) (-2.82901e-66,1.19825e-65) (1.18021e-66,1.82768e-66) (3.52604e-67,5.23873e-68) (4.01546e-68,-3.68127e-68) (-7.47986e-70,-7.76854e-69) (-9.19653e-70,-5.06808e-70) 
  (3.61395e-73,-3.807e-74) (-1.67724e-72,-2.95466e-72) (-1.75477e-71,2.45743e-71) (2.51938e-70,4.3082e-71) (-6.04207e-70,-1.96458e-69) (-1.10904e-68,1.10566e-68) (1.08223e-67,3.14584e-68) (-1.81769e-67,-7.41497e-67) (-3.43515e-66,3.42176e-66) (2.80203e-65,6.39425e-66) (-5.54798e-65,-1.48197e-64) (-4.62281e-64,6.59314e-64) (3.76934e-63,-2.36187e-65) (-9.63983e-63,-1.29891e-62) (-1.79833e-62,6.09462e-62) (2.12747e-61,-8.37623e-62) (-6.57939e-61,-3.63709e-61) (5.17577e-61,2.1651e-60) (2.88755e-60,-4.95834e-60) (-1.13822e-59,4.34124e-60) (1.90392e-59,4.2254e-60) (-1.53306e-59,-1.15739e-59) (6.40244e-60,-2.59929e-60) (-1.18832e-59,3.20287e-59) (1.38769e-59,-3.7715e-59) (3.07667e-59,1.26765e-59) (-8.21361e-59,1.75074e-59) (4.49081e-59,-6.25697e-59) (6.44013e-59,9.25733e-59) (-1.27427e-58,-9.41643e-60) (5.72824e-59,-1.22688e-58) (9.99562e-59,9.86122e-59) (-1.30008e-58,6.36921e-59) (-3.68557e-59,-1.14708e-58) (1.18177e-58,-2.08663e-59) (1.05548e-59,9.45716e-59) (-7.30961e-59,1.93204e-59) (-1.61301e-59,-6.58277e-59) (2.70854e-59,-3.22353e-59) (2.00727e-59,2.75781e-59) (6.34355e-60,2.83471e-59) (-4.03673e-60,2.22527e-60) (-9.0527e-60,-6.44639e-60) (-6.28955e-60,-1.91272e-60) (-1.72106e-60,6.98964e-61) (-5.30196e-63,1.04809e-61) (-9.5332e-62,-4.25913e-61) (-2.1414e-61,-3.04889e-61) (-1.0808e-61,-1.17654e-61) (-1.56689e-62,-4.99722e-62) (6.057e-63,-3.15033e-62) (1.8883e-63,-1.82511e-62) (-1.56215e-63,-7.77622e-63) (-1.58181e-63,-2.29446e-63) (-7.39815e-64,-3.87366e-64) (-2.1877e-64,1.64603e-65) (-3.93157e-65,3.31544e-65) (-1.97157e-66,1.07156e-65) (1.12476e-66,1.78181e-66) (3.66677e-67,7.8906e-68) (5.00396e-68,-3.63985e-68) (5.80775e-70,-9.49957e-69) (-1.03572e-69,-8.99714e-70) (-1.80003e-70,4.5665e-71) 
  (5.13344e-74,-4.583e-74) (-5.81329e-73,-2.63429e-73) (8.03861e-74,5.62474e-72) (4.2079e-71,-2.13953e-71) (-3.04587e-70,-2.20842e-70) (-3.86637e-70,2.81339e-69) (1.88495e-68,-7.36803e-69) (-1.06364e-67,-8.42558e-68) (-1.03977e-67,8.46115e-67) (4.51001e-66,-2.14973e-66) (-2.33165e-65,-1.39799e-65) (8.64896e-66,1.36432e-64) (4.91005e-64,-3.98918e-64) (-2.5996e-63,-6.80269e-64) (3.98332e-63,9.68412e-63) (1.84425e-62,-3.25916e-62) (-1.20201e-61,2.24626e-62) (2.88521e-61,2.11291e-61) (-1.73391e-61,-8.84747e-61) (-8.35557e-61,1.6484e-60) (2.40509e-60,-1.42538e-60) (-2.4027e-60,3.4286e-61) (-2.39707e-61,-1.23035e-60) (2.48347e-60,4.7281e-60) (-2.68462e-60,-4.39582e-60) (4.74055e-60,-3.66369e-60) (-5.86603e-60,1.12403e-59) (-4.25297e-60,-1.02448e-59) (1.75757e-59,5.88812e-61) (-1.20142e-59,1.43345e-59) (-1.00671e-59,-1.76662e-59) (2.07743e-59,-3.62724e-60) (-3.77581e-60,2.09041e-59) (-1.73176e-59,-5.11318e-60) (7.89478e-60,-1.58989e-59) (1.22243e-59,6.67316e-60) (-3.89266e-60,1.07798e-59) (-8.77845e-60,-3.78325e-60) (-1.72747e-60,-6.61735e-60) (4.38504e-60,4.89406e-62) (3.95063e-60,2.21668e-60) (3.26599e-61,7.52437e-61) (-1.44701e-60,2.72298e-61) (-9.16753e-61,4.68888e-61) (-1.61849e-61,3.01764e-61) (5.03295e-63,4.48562e-62) (-4.97492e-62,-2.61833e-62) (-5.52863e-62,-9.21048e-63) (-2.64782e-62,-6.66321e-64) (-8.56738e-63,-3.03258e-63) (-3.35363e-63,-3.67227e-63) (-1.98799e-63,-2.03771e-63) (-1.09103e-63,-6.23158e-64) (-4.46074e-64,-5.61259e-65) (-1.28358e-64,4.69996e-65) (-2.25912e-65,2.84612e-65) (-4.68793e-67,8.59114e-66) (1.07488e-66,1.49207e-66) (3.50534e-67,7.50826e-68) (5.39321e-68,-3.49807e-68) (1.73912e-69,-1.05359e-68) (-1.07591e-69,-1.25513e-69) (-2.39524e-70,1.11031e-71) (-1.75723e-71,2.75224e-71) 
  (2.76372e-75,-1.26156e-74) (-1.16315e-73,2.42912e-74) (6.29296e-73,8.26305e-73) (3.8256e-72,-7.74846e-72) (-6.8244e-71,1.33955e-72) (2.51625e-70,4.44096e-70) (1.85553e-69,-3.08747e-69) (-2.3903e-68,-1.95996e-70) (7.68599e-68,1.27132e-67) (3.79288e-67,-7.72843e-67) (-4.58998e-66,6.11981e-67) (1.54838e-65,1.70316e-65) (2.22892e-65,-1.02987e-64) (-4.04943e-64,1.80732e-64) (1.50308e-63,8.27687e-64) (-1.017e-63,-6.01595e-63) (-1.2627e-62,1.52084e-62) (5.68066e-62,-4.34071e-63) (-1.11357e-61,-8.50568e-62) (7.41375e-62,2.66352e-61) (1.08361e-61,-3.77571e-61) (-1.70478e-61,2.35699e-61) (-2.45007e-61,-6.85765e-62) (7.80726e-61,2.02e-61) (-6.29394e-61,-4.31199e-62) (-5.67314e-62,-1.0576e-60) (7.27519e-61,1.71271e-60) (-1.62117e-60,-2.39472e-61) (1.70951e-60,-2.08705e-60) (6.92319e-61,2.63052e-60) (-3.02372e-60,-3.08793e-61) (1.3696e-60,-2.83451e-60) (2.12844e-60,2.23342e-60) (-2.10623e-60,1.70294e-60) (-1.18537e-60,-2.30948e-60) (1.81734e-60,-9.0815e-61) (9.88362e-61,1.42097e-60) (-1.14258e-60,6.73233e-61) (-1.00665e-60,-4.16898e-61) (3.09356e-61,-4.54556e-61) (6.47334e-61,-2.16634e-61) (1.73652e-61,8.70615e-64) (-9.97366e-62,1.56327e-61) (-4.99504e-62,1.48082e-61) (1.35793e-62,5.85537e-62) (8.05086e-63,8.73045e-63) (-6.28369e-63,3.11561e-63) (-6.63877e-63,4.96326e-63) (-3.05661e-63,3.02639e-63) (-1.3238e-63,8.30748e-64) (-7.74023e-64,8.06521e-65) (-4.38314e-64,3.73512e-65) (-1.8644e-64,6.55967e-65) (-5.41779e-65,4.7418e-65) (-8.34408e-66,2.05902e-65) (9.23899e-67,5.90666e-66) (9.88059e-67,1.03417e-66) (3.0552e-67,4.26448e-68) (5.04645e-68,-3.36021e-68) (2.24254e-69,-1.07213e-68) (-1.05961e-69,-1.49474e-69) (-2.84341e-70,-2.57878e-71) (-2.87346e-71,3.0176e-71) (1.0662e-72,5.60855e-72) 
  (-9.64132e-76,-2.20042e-75) (-1.4646e-74,1.63199e-74) (1.82624e-73,5.27729e-74) (-2.88564e-73,-1.54127e-72) (-9.63442e-72,7.60702e-72) (8.37048e-71,3.55531e-71) (-7.43424e-71,-6.31164e-70) (-3.31121e-69,2.54153e-69) (2.40168e-68,9.04523e-69) (-3.12224e-68,-1.43715e-67) (-5.42004e-67,5.63871e-67) (3.79658e-66,6.08398e-67) (-7.75944e-66,-1.56022e-65) (-3.33134e-65,6.46528e-65) (2.7546e-64,-4.85298e-65) (-7.44274e-64,-6.51046e-64) (1.26757e-65,3.1742e-63) (6.33833e-63,-6.38366e-63) (-2.14677e-62,1.64787e-63) (3.4629e-62,2.14996e-62) (-2.49117e-62,-4.78887e-62) (6.53108e-63,3.16767e-62) (-3.78737e-62,3.04449e-62) (9.84064e-62,-6.4539e-62) (-4.16663e-62,6.22475e-62) (-1.48921e-61,-1.0213e-61) (2.55607e-61,7.29484e-62) (-1.58801e-61,1.92456e-61) (-9.03691e-62,-3.9622e-61) (3.70494e-61,1.3552e-61) (-2.99762e-61,3.37965e-61) (-2.21411e-61,-4.10888e-61) (4.40115e-61,-5.99318e-62) (2.77119e-62,4.04813e-61) (-3.7066e-61,-5.97573e-62) (4.1915e-62,-2.92904e-61) (2.59343e-61,5.12796e-63) (-1.41974e-62,1.81476e-61) (-1.47939e-61,8.24636e-62) (-3.09087e-62,-6.17373e-62) (4.01059e-62,-9.10721e-62) (1.96041e-62,-2.81596e-62) (5.85849e-63,2.10427e-62) (1.00406e-62,2.06867e-62) (8.32988e-63,5.76557e-63) (2.54721e-63,3.05761e-64) (-3.55807e-65,8.81229e-64) (-1.26103e-64,1.19933e-63) (1.35011e-65,6.85313e-64) (-3.40869e-65,2.628e-64) (-6.24696e-65,1.0592e-64) (-3.80985e-65,5.60871e-65) (-1.1207e-65,2.8786e-65) (-6.14933e-68,1.14477e-65) (1.56402e-66,3.22658e-66) (8.12875e-67,5.42118e-67) (2.3625e-67,-2.44239e-69) (4.02916e-68,-3.19672e-68) (1.85696e-69,-1.00223e-68) (-1.02434e-69,-1.54713e-69) (-3.07957e-70,-5.34911e-71) (-3.80243e-71,3.09492e-71) (3.28195e-74,7.19992e-72) (8.04932e-73,5.80616e-73) 
  (-3.82879e-76,-2.22821e-76) (-3.83865e-76,3.99322e-75) (3.22897e-74,-1.21252e-74) (-2.0826e-73,-1.90254e-73) (-5.45948e-73,2.11942e-72) (1.555e-71,-4.02734e-72) (-7.79246e-71,-7.92688e-71) (-1.8044e-70,6.99717e-70) (4.18957e-69,-1.32931e-69) (-1.92688e-68,-1.57902e-68) (-1.2199e-68,1.30465e-67) (5.54901e-67,-3.13725e-67) (-2.59536e-66,-1.20714e-66) (2.34721e-66,1.16267e-65) (2.9831e-65,-3.41765e-65) (-1.5931e-64,-4.97632e-66) (3.2796e-64,3.85447e-64) (9.11765e-65,-1.4041e-63) (-2.25583e-63,2.36586e-63) (5.80959e-63,-1.12304e-63) (-6.84623e-63,-2.33824e-63) (2.83674e-63,1.4618e-63) (-1.05555e-64,8.64195e-63) (2.5201e-63,-1.63942e-62) (5.23916e-63,7.63109e-63) (-2.84377e-62,8.34663e-63) (2.99686e-62,-2.17503e-62) (1.21546e-62,3.69402e-62) (-5.43531e-62,-2.55609e-62) (4.66667e-62,-3.31948e-62) (1.43897e-62,6.51127e-62) (-6.80657e-62,-9.26499e-63) (2.96085e-62,-5.61895e-62) (5.15564e-62,3.17492e-62) (-3.81998e-62,3.78103e-62) (-3.16009e-62,-2.9276e-62) (2.34646e-62,-3.04612e-62) (1.9639e-62,1.53801e-62) (-4.46296e-63,2.5249e-62) (-9.18173e-63,3.22929e-64) (-5.72991e-63,-1.28112e-62) (-1.73233e-63,-6.00542e-63) (2.14105e-63,9.31747e-64) (3.09332e-63,1.08332e-63) (1.6314e-63,-2.36819e-64) (4.0883e-64,-2.87686e-64) (1.14452e-64,5.00468e-65) (1.16661e-64,1.276e-64) (7.96197e-65,7.19827e-65) (2.97812e-65,3.26799e-65) (7.56045e-66,1.80703e-65) (3.06568e-66,9.97914e-66) (2.27658e-66,4.22623e-66) (1.35059e-66,1.20166e-66) (5.52132e-67,1.59538e-67) (1.54044e-67,-3.78215e-68) (2.61611e-68,-2.86241e-68) (7.58912e-70,-8.48894e-69) (-9.87853e-70,-1.38779e-69) (-3.06688e-70,-5.99911e-71) (-4.33944e-71,3.04602e-71) (-9.36344e-73,8.31884e-72) (8.62945e-73,8.86415e-73) (1.70009e-73,-2.31062e-74) 
  (-8.05354e-77,8.54888e-78) (3.75113e-76,6.23479e-76) (3.34439e-75,-5.22615e-75) (-5.00923e-74,-4.6789e-75) (1.50551e-73,3.56376e-73) (1.72689e-72,-2.22048e-72) (-1.91047e-71,-2.56171e-72) (4.96853e-71,1.13643e-70) (4.18838e-70,-6.17886e-70) (-4.18477e-69,-6.74929e-71) (1.19142e-68,1.82342e-68) (3.92555e-68,-9.73051e-68) (-4.54101e-67,1.10146e-67) (1.4761e-66,1.2344e-66) (2.72044e-67,-7.31635e-66) (-2.01861e-65,1.56518e-65) (7.90421e-65,1.28002e-65) (-1.32961e-64,-1.72625e-64) (-1.25204e-65,4.90001e-64) (4.98305e-64,-6.8249e-64) (-8.53701e-64,3.97554e-64) (2.08074e-64,-1.50173e-64) (1.07688e-63,9.70582e-64) (-1.443e-63,-1.73147e-63) (1.29554e-63,-4.15605e-64) (-1.89432e-63,4.2933e-63) (7.62753e-65,-5.04929e-63) (5.89369e-63,1.65407e-63) (-7.77436e-63,3.92631e-63) (-1.6091e-64,-8.34264e-63) (8.94296e-63,3.92517e-63) (-6.96461e-63,7.2195e-63) (-4.10699e-63,-8.05441e-63) (8.3032e-63,-3.41117e-63) (1.17403e-63,7.53607e-63) (-6.12531e-63,1.34942e-63) (-1.50793e-63,-5.41973e-63) (3.25218e-63,-1.16188e-63) (2.44785e-63,2.87813e-63) (-4.9548e-64,1.27288e-63) (-1.82232e-63,-5.80435e-64) (-9.67503e-64,-4.51935e-64) (1.7503e-64,-1.24367e-64) (4.06376e-64,-1.96823e-64) (1.60919e-64,-2.04108e-64) (1.90901e-65,-8.91473e-65) (1.53311e-65,-1.50906e-65) (2.44938e-65,-1.02455e-66) (1.6473e-65,-1.46182e-66) (7.25261e-66,-1.99738e-67) (3.03519e-66,7.86525e-67) (1.49674e-66,5.8663e-67) (7.26402e-67,1.52622e-67) (2.81414e-67,-3.52876e-68) (7.75769e-68,-4.8508e-68) (1.22532e-68,-2.24546e-68) (-5.11733e-70,-6.30341e-69) (-9.29032e-70,-1.05219e-69) (-2.79878e-70,-4.19317e-71) (-4.3146e-71,2.9605e-71) (-1.53865e-72,8.80833e-72) (8.77423e-73,1.1182e-72) (2.11276e-73,6.22995e-75) (1.84038e-74,-2.30485e-74) 
  (-1.08367e-77,9.90402e-78) (1.21038e-76,4.97414e-77) (-8.26044e-77,-1.10364e-75) (-7.55949e-75,4.69214e-75) (5.89153e-74,3.35696e-74) (1.70239e-75,-4.88435e-73) (-2.8626e-72,1.67055e-72) (1.85913e-71,1.00004e-71) (-9.08846e-72,-1.25397e-70) (-5.5359e-70,4.244e-70) (3.41058e-69,1.1325e-69) (-4.88237e-69,-1.64459e-68) (-4.64976e-68,5.99181e-68) (3.10556e-67,6.43692e-69) (-7.07358e-67,-9.39185e-67) (-8.74894e-67,3.9731e-66) (1.07181e-65,-6.55729e-66) (-3.27945e-65,-6.28266e-66) (4.74928e-65,5.48403e-65) (-1.43027e-65,-1.17725e-64) (-4.24464e-65,1.10467e-64) (-1.90958e-65,-1.43266e-65) (2.30619e-64,-2.321e-65) (-2.94387e-64,-3.37475e-66) (1.6363e-65,-2.37284e-64) (3.09601e-64,6.48555e-64) (-5.49693e-64,-3.99057e-64) (7.48708e-64,-6.0171e-64) (-2.36335e-64,1.21732e-63) (-1.02095e-63,-6.70639e-64) (1.22822e-63,-7.092e-64) (2.44681e-64,1.43232e-63) (-1.2724e-63,-1.75695e-64) (3.2268e-64,-1.27917e-63) (9.60876e-64,4.82024e-64) (-3.50143e-64,8.43067e-64) (-7.54958e-64,-2.97261e-64) (9.97131e-65,-4.78271e-64) (5.4189e-64,-6.20761e-66) (1.49059e-64,1.65072e-64) (-2.14756e-64,1.30392e-64) (-1.5984e-64,6.71771e-65) (-9.82921e-66,-1.56101e-65) (1.90652e-65,-5.67529e-65) (-3.95044e-66,-3.95934e-65) (-8.21597e-66,-1.35465e-65) (-1.08325e-66,-3.94311e-66) (2.0264e-66,-2.80712e-66) (1.5183e-66,-1.99939e-66) (7.44678e-67,-9.04098e-67) (3.97609e-67,-3.07174e-67) (2.13984e-67,-1.24976e-67) (8.98215e-68,-7.06667e-68) (2.46497e-68,-3.67169e-68) (2.44495e-69,-1.42616e-68) (-1.33832e-69,-3.87354e-69) (-8.05322e-70,-6.33797e-70) (-2.2962e-70,-7.68226e-72) (-3.70247e-71,2.85211e-71) (-1.50084e-72,8.5807e-72) (8.64771e-73,1.22502e-72) (2.38066e-73,3.02054e-74) (2.64787e-74,-2.42622e-74) (-4.53148e-76,-5.02199e-75) 
  (-5.08333e-79,2.5895e-78) (2.26066e-77,-5.79672e-78) (-1.29114e-76,-1.47143e-76) (-5.57344e-76,1.45739e-75) (1.1676e-74,-1.6035e-75) (-5.12346e-74,-6.66969e-74) (-2.09769e-73,5.24791e-73) (3.51091e-72,-6.09949e-73) (-1.41707e-71,-1.5506e-71) (-2.81968e-71,1.11867e-70) (5.52991e-70,-2.01964e-70) (-2.28336e-69,-1.59878e-69) (1.5684e-70,1.22444e-68) (3.95437e-68,-3.04477e-68) (-1.82479e-67,-4.46121e-68) (2.98258e-67,5.70382e-67) (5.92181e-67,-1.86262e-66) (-4.3417e-66,2.60095e-66) (1.05228e-65,1.21368e-66) (-1.25302e-65,-1.04729e-65) (5.60236e-66,1.30664e-65) (-3.7236e-66,5.143e-66) (2.13456e-65,-2.84456e-65) (-2.33752e-65,2.84621e-65) (-3.59625e-65,-2.40778e-65) (1.02881e-64,2.82185e-65) (-8.52954e-65,3.27193e-65) (-4.81989e-66,-1.48788e-64) (1.15493e-64,1.29679e-64) (-1.66451e-64,6.71276e-65) (2.26637e-65,-2.02896e-64) (1.86466e-64,9.38679e-65) (-1.23353e-64,1.34587e-64) (-1.20679e-64,-1.49143e-64) (1.32917e-64,-7.14377e-65) (7.05948e-65,1.12294e-64) (-9.83767e-65,6.01865e-65) (-5.17371e-65,-4.86034e-65) (4.7523e-65,-5.88824e-65) (3.65885e-65,-6.85214e-66) (-4.73725e-66,3.13471e-65) (-9.18286e-66,2.53661e-65) (-2.57856e-66,2.507e-66) (-3.52292e-66,-6.71642e-66) (-4.54087e-66,-3.79888e-66) (-2.55944e-66,-6.86053e-67) (-7.27553e-67,-2.67039e-67) (-1.51709e-67,-4.6863e-67) (-7.26488e-68,-3.69019e-67) (-3.02276e-68,-1.83685e-67) (9.09541e-70,-8.03153e-68) (5.29252e-69,-3.78797e-68) (4.67517e-70,-1.75297e-68) (-1.80665e-69,-6.61406e-69) (-1.42028e-69,-1.7756e-69) (-5.99775e-70,-2.56519e-70) (-1.62964e-70,2.59408e-71) (-2.6513e-71,2.63424e-71) (-8.24651e-73,7.62791e-72) (8.43338e-73,1.16938e-72) (2.46572e-73,4.14927e-74) (3.19553e-74,-2.45395e-74) (3.39482e-76,-6.05887e-75) (-6.47292e-76,-5.62154e-76) 
  (2.02222e-79,4.24755e-79) (2.58682e-78,-3.21666e-78) (-3.36307e-77,-6.94372e-78) (7.65709e-77,2.60349e-76) (1.42705e-75,-1.44588e-75) (-1.38929e-74,-3.64249e-75) (2.66499e-74,9.17912e-74) (3.99268e-73,-4.4342e-73) (-3.43637e-72,-5.63196e-73) (7.76411e-72,1.72752e-71) (5.0122e-71,-8.16436e-71) (-4.49498e-70,2.69806e-71) (1.24602e-69,1.5226e-69) (1.86629e-69,-7.76043e-69) (-2.68917e-68,1.29586e-68) (9.36609e-68,3.80826e-68) (-1.20167e-67,-2.76213e-67) (-2.23002e-67,7.24906e-67) (1.23193e-66,-8.985e-67) (-2.19868e-66,1.3066e-67) (1.48522e-66,6.08288e-67) (5.55893e-67,1.37513e-66) (-9.47698e-67,-5.172e-66) (1.13473e-66,4.25972e-66) (-7.13511e-66,2.72522e-66) (1.27619e-65,-8.57207e-66) (-2.18867e-66,1.23368e-65) (-1.8302e-65,-1.33686e-65) (2.38958e-65,-2.10634e-66) (-6.06791e-66,2.5688e-65) (-2.13915e-65,-1.97815e-65) (2.65464e-65,-1.3423e-65) (5.82796e-66,2.53447e-65) (-2.75582e-65,8.86566e-67) (2.38574e-66,-2.10242e-65) (1.9168e-65,1.1726e-66) (-1.52478e-66,1.60925e-65) (-1.02118e-65,2.64243e-66) (-2.14074e-66,-1.00632e-65) (2.56291e-66,-5.58132e-66) (2.64291e-66,2.77018e-66) (1.84568e-66,3.59629e-66) (3.0495e-67,8.20388e-67) (-8.75512e-67,-2.3417e-67) (-8.53018e-67,7.34668e-68) (-3.74756e-67,2.08941e-67) (-1.22021e-67,7.22311e-68) (-6.8701e-68,-2.03943e-68) (-4.83633e-68,-2.76665e-68) (-2.47706e-68,-1.537e-68) (-9.85841e-69,-8.12094e-69) (-4.08855e-69,-4.26634e-69) (-2.02318e-69,-1.76225e-69) (-9.55256e-70,-4.53439e-70) (-3.54668e-70,-1.74985e-71) (-9.37064e-71,4.31725e-71) (-1.46162e-71,2.19893e-71) (1.7279e-73,6.04017e-72) (8.07202e-73,9.57063e-73) (2.34709e-73,3.45996e-74) (3.36348e-74,-2.42367e-74) (8.92363e-76,-6.66754e-75) (-6.71601e-76,-7.67378e-76) (-1.44774e-76,7.59685e-78) 
  (7.35204e-80,3.89036e-80) (2.41367e-80,-7.23714e-79) (-5.39372e-78,2.57006e-78) (3.77626e-77,2.76667e-77) (4.24195e-77,-3.44722e-76) (-2.2373e-75,9.55476e-76) (1.30036e-74,9.3826e-75) (6.66648e-75,-9.8903e-74) (-5.01365e-73,2.77238e-73) (2.73904e-72,1.42515e-72) (-1.83513e-72,-1.53838e-71) (-5.39019e-71,4.82798e-71) (3.07671e-70,6.59613e-71) (-5.46867e-70,-1.14686e-69) (-1.96247e-69,4.28832e-69) (1.49555e-68,-4.97241e-69) (-4.16308e-68,-1.95046e-68) (4.75919e-68,1.01731e-67) (4.15125e-68,-2.12214e-67) (-1.98752e-67,2.11497e-67) (1.51675e-67,-6.35904e-68) (2.76708e-67,8.80738e-68) (-6.35155e-67,-4.0011e-67) (4.93976e-67,1.36156e-67) (-3.86049e-67,1.22995e-66) (2.45299e-67,-2.13929e-66) (1.36749e-66,1.14835e-66) (-3.26357e-66,8.80526e-67) (1.67946e-66,-2.8221e-66) (2.53191e-66,2.92873e-66) (-4.0504e-66,7.80227e-67) (7.03657e-67,-4.14556e-66) (3.45331e-66,1.37159e-66) (-2.26939e-66,3.18768e-66) (-2.24612e-66,-1.94716e-66) (1.7597e-66,-2.13244e-66) (1.66509e-66,1.49499e-66) (-5.19545e-67,1.49811e-66) (-1.2233e-66,-6.02339e-67) (-4.55545e-67,-8.71743e-67) (4.36933e-67,-7.42337e-68) (5.62773e-67,1.59126e-67) (1.72936e-67,5.04463e-68) (-8.22338e-68,5.65761e-68) (-7.68393e-68,9.24629e-68) (-1.89871e-68,6.47883e-68) (-4.60127e-69,2.45402e-68) (-8.27431e-69,6.93723e-69) (-7.68364e-69,2.82077e-69) (-4.30254e-69,1.32739e-69) (-1.97727e-69,3.94514e-70) (-9.09041e-70,8.61112e-71) (-4.03869e-70,6.80999e-71) (-1.48136e-70,6.62949e-71) (-3.8411e-71,3.9548e-71) (-4.81071e-72,1.54868e-71) (1.00376e-72,4.07674e-72) (7.27869e-73,6.42676e-73) (2.02727e-73,1.22075e-74) (3.0782e-74,-2.36417e-74) (1.0454e-75,-6.75451e-75) (-6.7735e-76,-8.88095e-76) (-1.6995e-76,-1.2797e-77) (-1.66023e-77,1.78571e-77) 
  (1.44145e-80,-2.24554e-81) (-7.23858e-80,-1.03137e-79) (-4.73109e-79,9.16201e-79) (8.00847e-78,-1.69424e-79) (-3.00184e-77,-5.06805e-77) (-1.98361e-76,3.57435e-76) (2.66701e-75,-1.02311e-76) (-9.20435e-75,-1.35038e-74) (-3.63222e-74,8.62412e-74) (4.91214e-73,-9.35311e-74) (-1.76503e-72,-1.75795e-72) (-1.95627e-72,1.14054e-71) (4.48096e-71,-2.24185e-71) (-1.81936e-70,-8.6096e-71) (1.95671e-70,7.1408e-70) (1.24914e-69,-2.09209e-69) (-6.65926e-69,1.97349e-69) (1.51694e-68,6.30733e-69) (-1.59449e-68,-2.56293e-68) (1.44217e-70,3.7232e-68) (5.01211e-69,-1.30667e-68) (4.42182e-68,-2.58615e-68) (-9.97415e-68,2.781e-68) (3.80319e-68,-4.89312e-68) (1.12209e-67,1.75744e-67) (-2.0262e-67,-2.12311e-67) (2.50407e-67,-8.90349e-68) (-2.01631e-67,4.50137e-67) (-1.85235e-67,-4.08386e-67) (5.62647e-67,-4.2933e-68) (-2.48123e-67,5.24109e-67) (-4.09359e-67,-4.24631e-67) (4.4392e-67,-2.93666e-67) (1.62407e-67,5.23577e-67) (-4.05539e-67,1.06774e-67) (-9.63053e-68,-3.83126e-67) (2.99972e-67,-6.43419e-68) (1.394e-67,1.93308e-67) (-1.57512e-67,7.99155e-68) (-1.49236e-67,-3.08263e-68) (1.55629e-68,-4.80801e-68) (6.97834e-68,-4.26239e-68) (2.76568e-68,-1.80802e-68) (-1.15975e-70,9.70738e-69) (1.7817e-69,1.62604e-68) (4.95012e-69,9.08572e-69) (2.55772e-69,3.38949e-69) (1.8582e-70,1.67862e-69) (-3.89606e-70,1.13146e-69) (-2.75584e-70,6.29015e-70) (-1.49366e-70,2.77935e-70) (-7.70187e-71,1.18062e-70) (-3.09012e-71,5.42081e-71) (-6.92899e-72,2.38127e-71) (6.88306e-73,8.48369e-72) (1.29991e-72,2.17463e-72) (5.8244e-73,3.17818e-73) (1.54348e-73,-1.50601e-74) (2.39281e-74,-2.23593e-74) (7.11008e-76,-6.2728e-75) (-6.70025e-76,-8.98063e-76) (-1.82796e-76,-2.443e-77) (-2.16064e-77,1.83213e-77) (9.03743e-80,4.0778e-78) 
  (1.77356e-81,-1.81574e-81) (-2.0699e-80,-6.68311e-81) (3.05385e-80,1.7388e-79) (1.06117e-78,-8.50194e-79) (-9.20991e-78,-3.65999e-78) (1.04683e-77,6.73424e-77) (3.36679e-76,-2.8457e-76) (-2.54912e-75,-8.08948e-76) (4.01659e-75,1.46387e-74) (5.27948e-74,-6.07475e-74) (-3.95806e-73,-4.57851e-74) (8.84964e-73,1.61578e-72) (3.31101e-72,-7.22103e-72) (-3.07734e-71,7.70245e-72) (9.51329e-71,6.54223e-71) (-6.59795e-71,-3.67579e-70) (-5.45044e-70,8.83671e-70) (2.23019e-69,-8.09187e-70) (-4.00097e-69,-1.07533e-69) (3.19573e-69,3.34508e-69) (-3.63574e-70,-5.56191e-70) (1.83995e-69,-8.22715e-69) (-6.036e-69,1.24012e-68) (-5.02925e-69,-7.28913e-69) (3.21184e-68,4.74532e-69) (-3.88532e-68,3.30132e-69) (8.86621e-69,-3.97906e-68) (3.13152e-68,6.30315e-68) (-6.06928e-68,-1.0236e-68) (4.39763e-68,-6.85957e-68) (3.8742e-68,7.1193e-68) (-8.14204e-68,1.08877e-68) (2.33088e-69,-7.62869e-68) (7.12658e-68,2.59055e-68) (-2.00088e-68,5.59932e-68) (-5.16767e-68,-2.14079e-68) (1.64864e-68,-3.84337e-68) (3.54928e-68,3.33148e-70) (-3.15402e-69,2.22887e-68) (-1.79594e-68,1.41251e-68) (-4.96963e-69,-3.80319e-69) (2.10878e-69,-1.08381e-68) (8.69038e-70,-5.54575e-69) (7.68675e-70,2.57603e-70) (1.71814e-69,1.29099e-69) (1.48605e-69,4.28183e-70) (6.9668e-70,7.18041e-71) (2.38709e-70,1.29517e-70) (9.46296e-71,1.47081e-70) (4.51633e-71,9.31987e-71) (1.83312e-71,4.53505e-71) (6.76781e-72,2.06306e-71) (3.4205e-72,8.85023e-72) (2.08846e-72,3.14422e-72) (1.05186e-72,7.75969e-73) (3.86415e-73,7.42917e-74) (9.85257e-74,-3.39945e-74) (1.4923e-74,-1.95815e-74) (3.10185e-77,-5.24942e-75) (-6.51242e-76,-7.86153e-76) (-1.81014e-76,-2.43223e-77) (-2.40109e-77,1.84516e-77) (-4.08276e-79,4.6652e-78) (4.84504e-79,4.75221e-79) 
  (5.67061e-83,-4.3445e-82) (-3.51772e-81,1.22585e-81) (2.20333e-80,2.03419e-80) (5.45092e-80,-2.22426e-79) (-1.59004e-78,4.57167e-79) (8.20653e-78,7.73131e-78) (1.47756e-77,-7.0743e-77) (-4.07103e-76,1.52038e-76) (1.96617e-75,1.45574e-75) (6.30802e-76,-1.2865e-74) (-5.39736e-74,3.33067e-74) (2.69245e-73,1.13141e-73) (-3.09703e-73,-1.21512e-72) (-2.94723e-72,4.0045e-72) (1.7779e-71,-1.8362e-72) (-4.43459e-71,-3.53575e-71) (2.76154e-71,1.50997e-70) (1.55488e-70,-3.00191e-70) (-4.92456e-70,2.63191e-70) (5.51641e-70,2.76771e-71) (7.21202e-71,6.26641e-71) (-7.39127e-70,-1.09045e-69) (7.10038e-70,1.62315e-69) (-1.46399e-69,3.21039e-70) (3.73563e-69,-3.14902e-69) (-2.72455e-69,4.2754e-69) (-4.31599e-69,-4.61043e-69) (9.5699e-69,2.21319e-69) (-5.83066e-69,6.25706e-69) (-3.95368e-69,-1.09372e-68) (1.11853e-68,1.45963e-69) (-5.44155e-69,9.98081e-69) (-8.67597e-69,-6.64825e-69) (8.68634e-69,-5.65549e-69) (4.93186e-69,6.8827e-69) (-6.73867e-69,4.00766e-69) (-3.03083e-69,-4.82313e-69) (3.19437e-69,-4.1134e-69) (2.17671e-69,1.86011e-69) (-1.3936e-70,3.31659e-69) (-7.72108e-70,5.39771e-70) (-8.68711e-70,-1.14412e-69) (-5.59529e-70,-7.0669e-70) (6.27328e-72,-1.0628e-70) (2.66099e-70,-5.24106e-71) (1.95847e-70,-1.11971e-70) (8.49367e-71,-7.36367e-71) (4.00326e-71,-1.88032e-71) (2.55914e-71,2.08722e-72) (1.49923e-71,3.80441e-72) (7.14934e-72,2.29932e-72) (3.11636e-72,1.18069e-72) (1.36928e-72,4.45478e-73) (5.68756e-73,6.43741e-74) (1.94864e-73,-4.3799e-74) (4.82181e-74,-3.69841e-74) (6.4109e-75,-1.49594e-74) (-6.68546e-76,-3.82732e-75) (-6.05425e-76,-5.77273e-76) (-1.63696e-76,-1.19022e-77) (-2.33058e-77,1.82524e-77) (-6.20296e-79,4.90555e-78) (4.92835e-79,5.91533e-79) (1.12314e-79,1.21707e-82) 
  (-3.69725e-83,-6.53012e-83) (-3.50563e-82,5.271e-82) (5.03225e-81,4.70928e-82) (-1.54376e-80,-3.50198e-80) (-1.61995e-79,2.21088e-79) (1.84303e-78,1.74967e-79) (-5.18929e-78,-1.0556e-77) (-3.66188e-77,5.98197e-77) (3.91737e-76,-1.08089e-77) (-1.18638e-75,-1.6726e-75) (-3.44293e-75,9.4429e-75) (4.43697e-74,-1.25494e-74) (-1.58192e-73,-1.17462e-73) (4.703e-74,7.73249e-73) (1.88768e-72,-1.99363e-72) (-8.52017e-72,4.35402e-73) (1.78212e-71,1.36322e-71) (-1.26437e-71,-4.57937e-71) (-2.35718e-71,6.99004e-71) (4.76037e-71,-4.05252e-71) (3.67169e-71,-8.45615e-72) (-1.94824e-70,-3.14612e-71) (2.11832e-70,5.67051e-71) (-8.06694e-71,2.52172e-70) (1.92151e-71,-7.12393e-70) (2.44513e-70,6.02545e-70) (-9.65189e-70,1.14666e-70) (1.06015e-69,-8.21926e-70) (2.85371e-70,1.1735e-69) (-1.55913e-69,-5.03117e-70) (1.07413e-69,-1.13849e-69) (6.69517e-70,1.41428e-69) (-1.49661e-69,4.3805e-70) (8.53573e-71,-1.3998e-69) (1.20824e-69,-9.45123e-72) (-1.14257e-70,1.08144e-69) (-7.79005e-70,-2.5865e-71) (-1.84472e-70,-7.27481e-70) (3.50649e-70,-1.25139e-70) (3.41473e-70,3.19654e-70) (2.9068e-71,1.58886e-70) (-1.79054e-70,-1.09141e-71) (-1.37888e-70,-1.10506e-71) (-2.51673e-71,-6.87011e-72) (1.57265e-71,-2.85998e-71) (7.68004e-72,-3.11902e-71) (7.16247e-73,-1.75879e-71) (1.58264e-72,-7.02336e-72) (2.51841e-72,-2.84929e-72) (1.85145e-72,-1.35104e-72) (9.65053e-73,-6.10608e-73) (4.40188e-73,-2.55813e-73) (1.83214e-73,-1.18174e-73) (6.26345e-74,-5.96558e-74) (1.4313e-74,-2.67891e-74) (6.53611e-76,-9.31048e-75) (-1.0551e-75,-2.29596e-75) (-5.12554e-76,-3.29911e-76) (-1.32327e-76,7.32177e-78) (-1.94528e-77,1.76047e-77) (-5.08067e-79,4.74379e-78) (4.9592e-79,6.31446e-79) (1.25354e-79,1.163e-80) (1.32041e-80,-1.29397e-80) 
  (-1.16985e-83,-5.07986e-84) (6.6642e-84,1.06538e-82) (7.16449e-82,-4.48652e-82) (-5.57107e-81,-3.04147e-81) (1.1807e-81,4.50506e-80) (2.54706e-79,-1.61844e-79) (-1.71063e-78,-8.29745e-79) (1.27971e-78,1.11751e-77) (4.80735e-77,-3.982e-77) (-3.11517e-76,-9.23558e-77) (4.98024e-76,1.50612e-75) (4.21036e-75,-5.90297e-75) (-3.07735e-74,1.45897e-75) (8.26432e-74,8.68961e-74) (1.83687e-74,-4.17865e-73) (-9.04044e-73,8.92741e-73) (3.22889e-72,-2.81764e-73) (-5.60227e-72,-3.44898e-72) (3.97625e-72,8.6613e-72) (7.69159e-73,-6.49497e-72) (4.25145e-72,-7.2949e-72) (-2.2554e-71,1.74227e-71) (2.02969e-71,-1.66407e-71) (2.72319e-71,3.64546e-71) (-7.35954e-71,-6.91102e-71) (8.20479e-71,1.58607e-71) (-7.61168e-71,1.25975e-70) (2.82737e-72,-1.7947e-70) (1.62438e-70,5.97161e-71) (-1.88235e-70,1.27976e-70) (-4.06079e-71,-2.12935e-70) (2.10859e-70,3.93514e-71) (-7.70689e-71,2.07221e-70) (-1.45268e-70,-1.19806e-70) (9.94963e-71,-1.40611e-70) (1.09757e-70,1.01208e-70) (-6.26281e-71,8.74921e-71) (-9.68463e-71,-4.32297e-71) (7.55496e-72,-5.02586e-71) (6.35568e-71,-7.1024e-72) (2.5989e-71,1.02282e-71) (-1.44002e-71,1.58093e-71) (-1.50543e-71,1.37879e-71) (-4.19343e-72,3.74321e-72) (-1.55906e-72,-3.37657e-72) (-2.44978e-72,-3.73085e-72) (-1.88819e-72,-1.9217e-72) (-7.1852e-73,-9.12359e-73) (-1.18519e-73,-5.57072e-73) (1.79043e-74,-3.37201e-73) (2.23372e-74,-1.70611e-73) (1.21896e-74,-7.63836e-74) (3.64902e-75,-3.27171e-74) (-8.53836e-76,-1.3e-74) (-1.66488e-75,-4.28611e-75) (-1.00128e-75,-1.01528e-75) (-3.72379e-76,-1.1618e-76) (-9.19845e-77,2.40668e-77) (-1.33981e-77,1.60085e-77) (-1.05542e-79,4.16871e-78) (4.89505e-79,5.87362e-79) (1.28847e-79,1.44571e-80) (1.57516e-80,-1.30773e-80) (5.26605e-83,-3.02628e-81) 
  (-2.0909e-84,5.0527e-85) (1.16776e-83,1.35179e-83) (4.91816e-83,-1.31414e-82) (-1.03207e-81,1.62671e-82) (4.6518e-81,5.69814e-81) (1.64938e-80,-4.59768e-80) (-2.9858e-79,6.3639e-80) (1.25671e-78,1.27912e-78) (2.11481e-78,-9.66371e-78) (-4.76516e-77,1.88935e-77) (2.08445e-76,1.36931e-76) (-6.66638e-77,-1.13345e-75) (-3.54688e-75,3.22175e-75) (1.83305e-74,1.95827e-75) (-3.94524e-74,-4.93345e-74) (-1.1218e-74,1.86934e-73) (3.1213e-73,-3.413e-73) (-8.7918e-73,1.77994e-73) (1.11251e-72,4.50198e-73) (-3.40441e-73,-4.90588e-73) (-4.2448e-73,-1.51564e-72) (-3.54606e-73,3.96421e-72) (-4.47088e-73,-3.06447e-72) (7.49071e-72,2.35449e-73) (-1.38489e-71,1.30331e-72) (7.32839e-72,-8.22138e-72) (7.39126e-72,2.05363e-71) (-1.83804e-71,-1.47805e-71) (2.04864e-71,-1.43719e-71) (-2.00366e-72,3.11253e-71) (-2.71445e-71,-1.27273e-71) (2.12064e-71,-2.02545e-71) (1.66796e-71,2.62313e-71) (-2.43147e-71,6.55677e-72) (-7.7249e-72,-2.32e-71) (1.99419e-71,-3.85299e-72) (5.31256e-72,1.4041e-71) (-1.30189e-71,6.80622e-72) (-5.86401e-72,-4.43027e-72) (4.69839e-72,-7.0652e-72) (3.93218e-72,-2.48259e-72) (5.10833e-73,2.36956e-72) (-1.16701e-74,2.90645e-72) (5.14507e-74,1.05798e-72) (-4.03395e-73,-3.42343e-74) (-5.97993e-73,-9.12221e-74) (-4.03441e-73,1.0771e-74) (-1.84674e-73,-5.66794e-75) (-7.8438e-74,-3.58485e-74) (-3.70084e-74,-3.29894e-74) (-1.74965e-74,-1.88311e-74) (-7.75448e-75,-8.73334e-75) (-3.46678e-75,-3.53966e-75) (-1.58187e-75,-1.15012e-75) (-6.54095e-76,-2.29237e-76) (-2.16382e-76,1.26297e-77) (-5.14549e-77,3.06455e-77) (-6.87821e-78,1.3045e-77) (4.03085e-79,3.24458e-78) (4.66485e-79,4.6557e-79) (1.21532e-79,8.8599e-81) (1.61469e-80,-1.31471e-80) (2.99909e-82,-3.29758e-81) (-3.40444e-82,-3.56407e-82) 
  (-2.28149e-85,2.78558e-85) (2.90306e-84,6.12112e-85) (-6.72911e-84,-2.21163e-83) (-1.17421e-82,1.23936e-82) (1.16128e-81,2.69439e-82) (-2.43531e-81,-7.46585e-81) (-3.13813e-80,3.72625e-80) (2.81808e-79,3.75412e-80) (-6.75557e-79,-1.40655e-78) (-4.05206e-78,6.96162e-78) (3.89009e-77,-3.54395e-78) (-1.19404e-76,-1.30681e-76) (-1.02753e-76,7.33822e-76) (2.31817e-75,-1.59322e-75) (-9.31166e-75,-1.63289e-75) (1.70716e-74,2.13145e-74) (-3.1986e-76,-6.51646e-74) (-6.96682e-74,9.80694e-74) (1.36656e-73,-5.31068e-74) (-3.73733e-74,-1.3408e-74) (-2.33574e-73,-1.27566e-73) (3.64705e-73,3.96055e-73) (-3.64726e-73,-1.10866e-73) (7.93959e-73,-8.79247e-73) (-1.08596e-72,1.51738e-72) (-4.86105e-73,-1.44148e-72) (2.97142e-72,1.08466e-72) (-2.96099e-72,7.59292e-73) (5.08e-74,-3.62338e-72) (3.1637e-72,2.78992e-72) (-3.62699e-72,1.99669e-72) (-5.62182e-73,-3.96448e-72) (4.3105e-72,3.80135e-73) (-1.13385e-72,3.17418e-72) (-3.27003e-72,-1.08776e-72) (1.16202e-72,-2.48519e-72) (2.05758e-72,4.85708e-73) (-3.64592e-73,1.96182e-72) (-1.02324e-72,4.20797e-73) (-3.24692e-73,-1.04297e-72) (8.22077e-74,-7.36092e-73) (2.52837e-73,7.81046e-74) (2.94566e-73,2.70217e-73) (1.4357e-73,1.13297e-73) (-1.81633e-74,4.25169e-74) (-6.07263e-74,5.20028e-74) (-3.89564e-74,4.46224e-74) (-1.94881e-74,2.13774e-74) (-1.15697e-74,6.28547e-75) (-7.15868e-75,1.26924e-75) (-3.80369e-75,2.28858e-76) (-1.75058e-75,6.7797e-77) (-7.39879e-76,6.63063e-77) (-2.83612e-76,7.20457e-77) (-8.98768e-77,5.24118e-77) (-2.00969e-77,2.59035e-77) (-1.74593e-78,8.97742e-78) (7.72078e-79,2.13957e-78) (4.12963e-79,2.97906e-79) (1.03538e-79,-3.0086e-81) (1.43626e-80,-1.29116e-80) (3.00812e-82,-3.31218e-81) (-3.42462e-82,-4.07988e-82) (-7.98058e-83,-2.12283e-84) 
  (-2.28709e-87,5.97755e-86) (4.41884e-85,-2.09675e-85) (-3.07304e-84,-2.20247e-84) (-2.83426e-84,2.75533e-83) (1.74432e-82,-7.99466e-83) (-1.03789e-81,-7.04584e-82) (-3.07864e-82,7.72282e-81) (3.87239e-80,-2.2623e-80) (-2.19622e-79,-1.08781e-79) (1.76108e-79,1.24873e-78) (4.39512e-78,-4.22251e-78) (-2.71788e-77,-3.97247e-78) (6.04497e-77,9.65021e-77) (1.07667e-76,-4.11982e-76) (-1.19253e-75,7.36173e-76) (3.88998e-75,6.15481e-76) (-6.19704e-75,-6.6104e-75) (2.16719e-75,1.56969e-74) (7.46154e-75,-1.55508e-74) (-5.10283e-76,-1.68583e-75) (-4.03371e-74,1.24391e-74) (7.05958e-74,-1.49189e-75) (-3.32821e-74,4.13176e-74) (-2.09179e-74,-1.79295e-73) (5.97312e-74,2.36549e-73) (-2.16331e-73,-4.49456e-74) (3.89302e-73,-2.21248e-73) (-1.41524e-73,3.67266e-73) (-4.12789e-73,-3.19302e-73) (5.5317e-73,-1.09449e-73) (-7.35736e-74,5.65805e-73) (-4.85119e-73,-2.52218e-73) (4.04458e-73,-4.37354e-73) (2.67608e-73,3.66449e-73) (-3.97051e-73,2.71585e-73) (-1.81278e-73,-3.21382e-73) (2.21947e-73,-2.00828e-73) (1.77523e-73,1.98237e-73) (-3.15702e-74,1.65736e-73) (-1.2809e-73,-4.74373e-74) (-7.82319e-74,-8.17866e-74) (1.81235e-74,-2.42139e-74) (5.28183e-74,-5.3916e-75) (2.92485e-74,-5.0771e-75) (5.58549e-75,3.9138e-75) (2.66079e-76,1.03108e-74) (9.88083e-76,8.46745e-75) (5.17278e-76,4.42302e-75) (-3.1381e-76,1.99361e-75) (-4.97983e-76,9.43699e-76) (-3.28064e-76,4.55267e-76) (-1.57721e-76,2.0799e-76) (-6.23463e-77,9.17103e-77) (-1.8741e-77,3.93978e-77) (-2.72696e-78,1.5314e-77) (9.55193e-79,4.84224e-78) (8.42364e-79,1.10484e-78) (3.22577e-79,1.33002e-79) (7.73058e-80,-1.56008e-80) (1.0754e-80,-1.21015e-80) (9.66921e-83,-3.0427e-81) (-3.43624e-82,-4.01343e-82) (-8.49506e-83,-6.95569e-84) (-9.35087e-84,8.83326e-84) 
  (5.65253e-87,8.08429e-87) (3.67263e-86,-7.11198e-86) (-6.13615e-85,1.94635e-86) (2.34445e-84,3.79738e-84) (1.42733e-83,-2.71603e-83) (-1.988e-82,1.23307e-83) (7.08176e-82,9.93031e-82) (2.62097e-81,-6.53682e-81) (-3.75558e-80,7.75478e-81) (1.4235e-79,1.35799e-79) (1.20802e-79,-9.39454e-79) (-3.62745e-78,2.1957e-78) (1.65646e-77,5.26765e-78) (-2.84826e-77,-5.72295e-77) (-5.82871e-77,1.97292e-76) (4.68232e-76,-3.09963e-76) (-1.23977e-75,-8.33037e-77) (1.59441e-75,1.28298e-75) (-5.7001e-76,-1.84471e-75) (-1.6355e-76,-9.07959e-76) (-2.88751e-75,5.69314e-75) (5.65773e-75,-6.98259e-75) (3.70326e-75,7.5103e-75) (-2.1762e-74,-1.53259e-74) (2.82375e-74,1.31612e-74) (-2.31162e-74,2.37501e-74) (1.17755e-74,-6.07812e-74) (2.91469e-74,4.1729e-74) (-7.20086e-74,1.85413e-74) (3.24499e-74,-6.72816e-74) (5.64906e-74,5.43368e-74) (-6.65996e-74,3.39023e-74) (-1.32515e-74,-7.9953e-74) (6.16512e-74,-2.41763e-75) (-3.62772e-75,6.62917e-74) (-4.93565e-74,-4.82367e-75) (-5.08728e-75,-4.20826e-74) (3.4796e-74,-3.05323e-75) (1.76967e-74,1.84062e-74) (-1.37654e-74,9.39343e-75) (-1.66295e-74,9.35745e-76) (-2.69854e-75,-3.31559e-75) (3.88053e-75,-5.5847e-75) (2.4531e-75,-3.88381e-75) (1.02699e-75,-6.96836e-76) (1.0642e-75,7.54412e-76) (9.86045e-76,6.90764e-76) (5.55457e-76,3.81739e-76) (2.10826e-76,2.26105e-76) (6.51856e-77,1.42769e-76) (2.16324e-77,7.92887e-77) (9.00188e-78,3.7572e-77) (4.65972e-78,1.58041e-77) (2.72752e-78,5.87873e-78) (1.47763e-78,1.78375e-78) (6.41971e-79,3.67245e-79) (2.09411e-79,1.55224e-80) (4.80706e-80,-2.2878e-80) (6.30562e-81,-1.03827e-80) (-2.27409e-82,-2.50614e-81) (-3.34532e-82,-3.40364e-82) (-8.33243e-83,-5.20086e-84) (-1.02812e-83,8.85238e-84) (-5.88035e-86,2.06107e-84) 
  (1.53694e-87,4.95435e-88) (-2.25794e-87,-1.2808e-86) (-7.66587e-86,6.26417e-86) (6.6786e-85,2.53297e-85) (-8.37758e-85,-4.80338e-84) (-2.36539e-83,2.07259e-83) (1.834e-82,5.52506e-83) (-3.03632e-82,-1.05877e-81) (-3.86459e-81,4.56232e-81) (3.04578e-80,2.77312e-81) (-7.70111e-80,-1.24714e-79) (-2.12558e-79,6.15219e-79) (2.42628e-78,-1.02577e-78) (-8.80847e-78,-3.59329e-78) (1.29173e-77,2.69576e-77) (1.89176e-77,-7.68283e-77) (-1.29983e-76,1.0633e-76) (2.57711e-76,-2.04336e-77) (-1.7284e-76,-1.02972e-76) (-1.71176e-76,-1.49425e-76) (3.07855e-76,8.76294e-76) (-2.41217e-76,-1.08637e-75) (1.38083e-75,1.06894e-76) (-3.71526e-75,8.42334e-76) (3.46494e-75,-1.79333e-75) (9.41202e-76,4.92415e-75) (-5.20004e-75,-6.54935e-75) (6.69315e-75,-2.52478e-76) (-4.2684e-75,9.53404e-75) (-4.59974e-75,-8.69781e-75) (1.05767e-74,-1.74948e-75) (-1.54347e-75,1.01101e-74) (-9.58462e-75,-5.17819e-75) (4.45781e-75,-7.2244e-75) (6.85508e-75,5.90775e-75) (-4.31027e-75,5.11055e-75) (-5.22709e-75,-2.89598e-75) (2.31583e-75,-3.89653e-75) (3.76576e-75,-4.58919e-76) (7.56774e-77,2.01001e-75) (-1.44006e-75,1.87932e-75) (-6.94119e-76,2.28649e-76) (-2.33519e-76,-8.05191e-76) (-1.84435e-76,-6.57756e-76) (-1.34511e-77,-2.27823e-76) (1.5296e-76,-5.84466e-77) (1.6202e-76,-4.04511e-77) (9.72076e-77,-2.47667e-77) (4.70011e-77,-3.5935e-78) (2.25529e-77,5.20929e-78) (1.0997e-77,4.76841e-78) (5.11572e-78,2.4732e-78) (2.24291e-78,9.49836e-79) (9.2721e-79,2.44369e-79) (3.43525e-79,3.34966e-81) (1.0407e-79,-3.66359e-80) (2.26006e-80,-2.20581e-80) (2.30638e-81,-7.74406e-81) (-5.17728e-82,-1.78753e-81) (-3.06961e-82,-2.38981e-82) (-7.44015e-83,1.20772e-84) (-9.69189e-84,8.84543e-84) (-1.40983e-85,2.14361e-84) (2.26184e-85,2.38671e-85) 
  (2.47687e-88,-8.68367e-89) (-1.54245e-87,-1.42295e-87) (-3.65474e-87,1.54306e-86) (1.0879e-85,-3.27172e-86) (-5.67687e-85,-5.2078e-85) (-9.54625e-85,4.84716e-84) (2.79694e-83,-1.07078e-83) (-1.38617e-82,-1.01202e-82) (-3.4348e-83,9.28511e-82) (3.95454e-81,-2.60821e-81) (-2.13401e-80,-7.37094e-81) (3.55159e-80,9.27415e-80) (1.75305e-79,-3.5526e-79) (-1.32331e-78,4.65766e-79) (3.98133e-78,1.61977e-78) (-5.33749e-78,-9.63357e-78) (-2.90712e-78,2.21576e-77) (2.13461e-77,-2.36172e-77) (-1.83917e-77,2.99568e-78) (-4.37415e-77,1.26487e-78) (1.19413e-76,5.31896e-77) (-1.23971e-76,-5.3665e-77) (1.44824e-76,-1.74179e-76) (-2.59923e-76,4.62326e-76) (6.95599e-77,-4.78383e-76) (6.74079e-76,3.32677e-76) (-1.10338e-75,-3.70304e-77) (4.54264e-76,-7.838e-76) (6.514e-76,1.28862e-75) (-1.28191e-75,-1.78353e-76) (6.74313e-76,-1.29281e-75) (9.98443e-76,9.82581e-76) (-1.32208e-75,5.89087e-76) (-4.80597e-76,-1.07821e-75) (1.19252e-75,-2.46531e-76) (2.4351e-76,8.73505e-76) (-7.59412e-76,3.48123e-76) (-2.46238e-76,-5.31341e-76) (2.83588e-76,-4.72154e-76) (2.22546e-76,1.09044e-76) (6.78198e-77,3.18552e-76) (-2.59037e-77,1.25447e-76) (-9.32606e-77,-3.451e-77) (-8.80927e-77,-4.31507e-77) (-3.35426e-77,-2.15225e-77) (3.37696e-78,-2.06697e-77) (1.00143e-77,-2.0462e-77) (6.62708e-78,-1.31087e-77) (4.06419e-78,-5.86184e-78) (2.64379e-78,-2.17159e-78) (1.53742e-78,-8.20832e-79) (7.52704e-79,-3.51531e-79) (3.17214e-79,-1.66358e-79) (1.14883e-79,-8.22364e-80) (3.30888e-80,-3.84763e-80) (5.96595e-81,-1.52615e-80) (-2.4311e-82,-4.72042e-81) (-6.37212e-82,-1.04051e-81) (-2.54198e-82,-1.25736e-82) (-5.90608e-83,9.47493e-84) (-7.80258e-84,8.50193e-84) (-5.58058e-86,2.05052e-84) (2.25713e-85,2.52084e-85) (5.21556e-86,1.22755e-87) 
  (2.3374e-89,-3.53368e-89) (-3.34889e-88,-3.1597e-89) (1.02952e-87,2.30454e-87) (1.0505e-86,-1.45697e-86) (-1.20609e-85,-1.05582e-86) (3.44111e-85,6.91582e-85) (2.42663e-84,-3.98367e-84) (-2.66414e-83,8.26007e-85) (8.4888e-83,1.16215e-82) (2.23349e-82,-6.95963e-82) (-3.2421e-81,1.20834e-81) (1.31947e-80,7.2433e-81) (-1.51048e-80,-5.71351e-80) (-9.87341e-80,1.79582e-79) (5.73379e-79,-2.12195e-79) (-1.43922e-78,-4.68743e-79) (1.71374e-78,2.37017e-78) (-7.90894e-80,-3.80173e-78) (-1.01506e-78,9.0742e-79) (-5.23283e-78,5.3677e-78) (1.64232e-77,-7.01431e-78) (-1.35792e-77,9.17505e-78) (-7.46317e-78,-3.51353e-77) (2.30313e-77,6.81557e-77) (-4.50704e-77,-3.99511e-77) (1.00317e-76,-4.68338e-77) (-9.50634e-77,1.06227e-76) (-5.76599e-77,-1.12159e-76) (1.9149e-76,4.26184e-77) (-1.16925e-76,1.24513e-76) (-8.43721e-77,-1.78058e-76) (1.89319e-76,-3.10588e-77) (-4.35628e-77,1.85214e-76) (-1.62286e-76,-3.12957e-77) (7.00126e-77,-1.45889e-76) (1.17424e-76,3.96311e-77) (-2.41775e-77,1.12964e-76) (-7.53032e-77,-1.0789e-77) (-2.73558e-77,-7.30669e-77) (2.54853e-77,-2.03432e-77) (3.83159e-77,2.03827e-77) (1.4719e-77,1.57038e-77) (-9.09936e-78,6.95015e-78) (-1.25874e-77,5.25489e-78) (-6.25091e-78,2.11725e-78) (-2.27313e-78,-1.69083e-78) (-1.28989e-78,-2.77865e-78) (-8.02806e-79,-1.95916e-78) (-2.90826e-79,-1.02857e-78) (-1.45081e-80,-5.05982e-79) (4.46028e-80,-2.48934e-79) (2.92195e-80,-1.17215e-79) (1.06001e-80,-5.13114e-80) (1.45483e-81,-2.06754e-80) (-1.1966e-81,-7.36904e-81) (-1.13703e-81,-2.13966e-81) (-5.52463e-82,-4.3649e-82) (-1.80335e-82,-3.2925e-83) (-4.00523e-83,1.5626e-83) (-5.08482e-84,7.60544e-84) (1.26807e-85,1.77548e-84) (2.23948e-85,2.27122e-85) (5.29655e-86,2.27468e-87) (5.92991e-87,-5.71332e-87) 
  (-4.40288e-91,-6.78012e-90) (-4.54899e-89,2.83104e-89) (3.50765e-88,1.9096e-88) (-8.05186e-89,-2.82338e-87) (-1.59731e-86,1.01687e-86) (1.08129e-85,5.26916e-86) (-8.02838e-86,-7.19512e-85) (-3.17225e-84,2.63907e-84) (2.14151e-83,5.9148e-84) (-4.06598e-83,-1.04683e-82) (-2.62085e-82,4.57542e-82) (2.2176e-81,-4.62553e-82) (-7.25812e-81,-4.87204e-81) (6.77972e-81,2.88605e-80) (3.9132e-80,-7.65811e-80) (-1.85941e-79,8.69939e-80) (3.69397e-79,6.97894e-80) (-3.05531e-79,-3.12771e-79) (-7.20051e-80,2.9937e-80) (1.00588e-80,1.19515e-78) (7.75754e-79,-2.2434e-78) (1.80968e-79,2.05234e-78) (-4.85805e-78,-2.58937e-78) (8.76221e-78,3.7179e-78) (-7.3724e-78,2.29362e-78) (4.08245e-78,-1.54217e-77) (2.83152e-78,1.78078e-77) (-1.77976e-77,-2.09704e-78) (2.06377e-77,-1.61217e-77) (4.65918e-78,2.22223e-77) (-2.5878e-77,-5.42162e-78) (1.19717e-77,-2.33404e-77) (1.5947e-77,1.89871e-77) (-1.68469e-77,1.59202e-77) (-9.81528e-78,-1.88594e-77) (1.36322e-77,-1.02461e-77) (1.0372e-77,1.18929e-77) (-6.45946e-78,7.69119e-78) (-1.0247e-77,-3.35345e-78) (-1.06427e-78,-4.55921e-78) (5.16677e-78,-2.17462e-78) (3.42539e-78,-3.1662e-79) (2.59247e-79,1.30558e-78) (-5.63068e-79,1.75183e-78) (-3.76004e-79,9.74547e-79) (-3.70961e-79,1.83537e-79) (-3.9745e-79,-9.05067e-80) (-2.8546e-79,-9.43491e-80) (-1.44784e-79,-6.42859e-80) (-6.02662e-80,-4.4356e-80) (-2.4398e-80,-2.73503e-80) (-1.055e-80,-1.39405e-80) (-4.80101e-81,-5.9224e-81) (-2.19124e-81,-2.08827e-81) (-9.39359e-82,-5.60145e-82) (-3.48137e-82,-7.78053e-83) (-1.02635e-82,1.90594e-83) (-2.16201e-83,1.68428e-83) (-2.31908e-84,6.05554e-84) (3.23951e-85,1.35378e-84) (2.11712e-85,1.72552e-85) (4.93285e-86,-7.37349e-88) (6.00887e-87,-5.67046e-87) (1.55684e-89,-1.2928e-87) 
  (-7.09093e-91,-8.1848e-91) (-3.0195e-90,7.92911e-90) (6.21146e-89,-9.56657e-90) (-2.78184e-88,-3.43417e-88) (-1.0122e-87,2.76941e-87) (1.82818e-86,-3.74306e-87) (-7.79745e-86,-8.04151e-86) (-1.34081e-85,6.22616e-85) (3.14218e-84,-1.3439e-84) (-1.49458e-83,-8.46084e-84) (1.41678e-83,7.86042e-83) (2.05559e-82,-2.68781e-82) (-1.27017e-81,1.71432e-82) (3.49677e-81,2.40808e-81) (-3.24184e-81,-1.1511e-80) (-1.01429e-80,2.55147e-80) (3.98042e-80,-2.5661e-80) (-4.77256e-80,-2.4215e-81) (-2.38777e-80,8.99291e-82) (1.29682e-79,1.2644e-79) (-1.51933e-79,-2.67503e-79) (2.58446e-79,1.05271e-79) (-7.63629e-79,2.90332e-79) (1.10642e-78,-5.3665e-79) (-2.33452e-79,1.01185e-78) (-1.2737e-78,-1.85001e-78) (1.96053e-78,1.0863e-78) (-1.72503e-78,1.90111e-78) (8.05701e-80,-3.43488e-78) (2.80266e-78,1.19434e-78) (-2.65944e-78,2.3105e-78) (-1.56902e-78,-3.21187e-78) (3.20557e-78,-2.21259e-79) (3.90137e-79,3.21623e-78) (-2.7364e-78,-4.20171e-79) (-8.71657e-80,-2.35476e-78) (2.12269e-78,-1.6166e-79) (4.34143e-79,1.28702e-78) (-1.21403e-78,8.00762e-79) (-6.87306e-79,-1.88344e-79) (1.81543e-79,-6.78782e-79) (2.93035e-79,-4.36199e-79) (1.68639e-79,2.67722e-80) (1.3063e-79,2.02766e-79) (7.61207e-80,1.39748e-79) (-3.29213e-81,6.40098e-80) (-4.08037e-80,3.53675e-80) (-3.58641e-80,2.2043e-80) (-2.08203e-80,1.02399e-80) (-1.06362e-80,2.92563e-81) (-5.29567e-81,3.43531e-82) (-2.51857e-81,-7.11583e-83) (-1.10368e-81,-3.87103e-84) (-4.36923e-82,5.22033e-83) (-1.50661e-82,5.24965e-83) (-4.182e-83,3.13898e-83) (-7.83278e-84,1.32654e-83) (-2.64552e-85,4.06874e-84) (4.39866e-85,8.68027e-85) (1.83907e-85,1.02863e-85) (4.13207e-86,-5.55494e-87) (5.15532e-87,-5.57157e-87) (1.68848e-89,-1.28069e-87) (-1.42243e-88,-1.43316e-88) 
  (-1.6791e-91,-3.54909e-92) (3.76486e-91,1.28215e-90) (6.83294e-90,-7.08069e-90) (-6.68902e-89,-1.62682e-89) (1.36231e-88,4.36607e-88) (1.88828e-87,-2.18192e-87) (-1.71077e-86,-2.42446e-87) (4.30748e-86,8.8016e-86) (2.46137e-85,-4.62199e-85) (-2.57334e-84,4.53821e-85) (9.27566e-84,7.64354e-84) (-3.20048e-84,-5.0042e-83) (-1.20995e-82,1.41537e-82) (5.96118e-82,-8.2387e-83) (-1.40392e-81,-8.54027e-82) (1.3378e-81,3.36225e-81) (1.37404e-81,-5.66765e-81) (-3.76859e-81,3.05227e-81) (-4.78113e-81,3.33561e-81) (2.63781e-80,-6.45762e-82) (-3.8316e-80,-7.15657e-81) (3.16304e-80,-2.58602e-80) (-4.20765e-80,1.09929e-79) (3.88229e-80,-1.50422e-79) (1.0517e-79,1.02119e-79) (-3.06911e-79,-3.52856e-80) (2.50724e-79,-1.14186e-79) (6.84006e-80,3.6011e-79) (-3.37938e-79,-2.87081e-79) (3.50766e-79,-2.16879e-79) (3.16815e-80,4.65252e-79) (-4.75596e-79,-9.32003e-80) (2.16512e-79,-3.55045e-79) (3.88385e-79,2.26087e-79) (-2.49791e-79,2.57391e-79) (-2.72624e-79,-1.78221e-79) (1.50782e-79,-2.40484e-79) (1.83419e-79,4.21347e-80) (-1.52237e-80,1.9109e-79) (-8.09032e-80,7.4549e-80) (-5.43081e-80,-6.64057e-80) (-2.17529e-80,-7.40215e-80) (1.2601e-80,-2.228e-80) (3.06772e-80,2.72644e-81) (2.29578e-80,4.81741e-81) (8.27575e-81,5.8571e-81) (7.75811e-82,7.14174e-81) (-8.1102e-82,5.76288e-81) (-7.95865e-82,3.26175e-81) (-6.36503e-82,1.48828e-81) (-4.32534e-82,6.34195e-82) (-2.33614e-82,2.76302e-82) (-1.00812e-82,1.22946e-82) (-3.44088e-83,5.35727e-83) (-8.20023e-84,2.16754e-83) (-4.721e-85,7.61699e-84) (7.16006e-85,2.14669e-84) (4.24841e-85,4.28845e-85) (1.4022e-85,3.81109e-86) (3.01503e-86,-9.91288e-87) (3.66863e-87,-5.16134e-87) (-7.48785e-89,-1.15961e-87) (-1.40302e-88,-1.39041e-88) (-3.13692e-89,2.00665e-91) 
  (-2.44847e-92,1.15084e-92) (1.68355e-91,1.24523e-91) (1.8109e-91,-1.52279e-90) (-9.78583e-90,4.27487e-90) (5.77048e-89,4.08395e-89) (2.55191e-89,-4.44098e-88) (-2.30496e-87,1.32276e-87) (1.35605e-86,6.47327e-87) (-1.52517e-86,-7.84217e-86) (-2.55247e-85,3.01887e-85) (1.7957e-84,-3.36301e-86) (-5.20899e-84,-5.21307e-84) (6.92914e-85,2.6789e-83) (5.37047e-83,-6.51e-83) (-2.18322e-82,4.56205e-83) (4.26155e-82,1.96932e-82) (-3.49252e-82,-6.05819e-82) (-8.58335e-83,4.26112e-82) (-2.78364e-82,1.08355e-81) (2.51274e-81,-2.74414e-81) (-3.67374e-81,3.16649e-81) (-7.96732e-82,-6.18593e-81) (7.47978e-81,1.47128e-80) (-1.13876e-80,-1.55093e-80) (2.08077e-80,-4.63068e-81) (-3.08084e-80,2.78358e-80) (6.01033e-81,-3.33198e-80) (4.59001e-80,2.39425e-80) (-5.53166e-80,1.09688e-80) (3.89099e-81,-5.60268e-80) (5.1476e-80,3.34452e-80) (-4.88569e-80,4.32797e-80) (-2.20197e-80,-4.93474e-80) (5.71055e-80,-2.32748e-80) (9.14449e-81,4.55758e-80) (-4.18636e-80,1.61144e-80) (-1.40086e-80,-3.47578e-80) (1.88795e-80,-1.86303e-80) (1.84838e-80,1.64464e-80) (2.30284e-81,1.65926e-80) (-1.02479e-80,1.16009e-81) (-1.00319e-80,-4.34836e-81) (-2.35813e-81,-3.46101e-81) (2.5198e-81,-2.9135e-81) (2.65016e-81,-2.06352e-81) (1.50049e-81,-5.39362e-82) (8.6257e-82,4.4294e-82) (5.43276e-82,5.81423e-82) (2.85209e-82,3.86093e-82) (1.11087e-82,2.08272e-82) (3.36322e-83,1.05667e-82) (1.016e-83,5.07959e-83) (4.58066e-84,2.23325e-83) (2.80483e-84,8.73059e-84) (1.64501e-84,2.92031e-84) (7.98917e-85,7.69226e-85) (3.05797e-85,1.26431e-85) (8.87952e-86,-5.07958e-87) (1.81458e-86,-1.16974e-86) (1.95655e-87,-4.33532e-87) (-1.92898e-88,-9.37342e-88) (-1.36129e-88,-1.1314e-88) (-3.03023e-89,7.31833e-91) (-3.36424e-90,3.49146e-90) 
  (-1.97893e-93,3.75412e-93) (3.26576e-92,-3.28522e-94) (-1.2021e-91,-2.05364e-91) (-8.04687e-91,1.44081e-90) (1.08844e-89,-3.97472e-91) (-3.85867e-89,-5.64449e-89) (-1.53292e-88,3.77575e-88) (2.23603e-87,-5.20071e-88) (-9.33345e-87,-7.74776e-87) (-1.61911e-88,5.94437e-86) (1.98263e-85,-1.7791e-85) (-1.0718e-84,-6.48334e-86) (2.63877e-84,2.76123e-84) (-6.67698e-85,-1.16873e-83) (-1.71116e-83,2.45027e-83) (5.66741e-83,-1.93138e-83) (-7.78514e-83,-2.30072e-83) (9.92815e-84,2.85225e-83) (9.12791e-83,1.67281e-82) (-3.66901e-83,-5.0882e-82) (4.17125e-83,5.9612e-82) (-8.449e-82,-4.48337e-82) (2.17687e-81,5.95178e-82) (-2.34727e-81,-6.00907e-83) (1.22648e-81,-2.87085e-81) (6.98065e-83,5.45457e-81) (-3.08566e-81,-2.89056e-81) (6.61854e-81,-2.83334e-81) (-3.15386e-81,6.35012e-81) (-5.84274e-81,-4.95754e-81) (7.54743e-81,-2.79546e-81) (6.07349e-82,8.69939e-81) (-6.98168e-81,-1.22312e-81) (2.26874e-81,-8.03852e-81) (5.61043e-81,2.30427e-81) (-1.59928e-81,5.92224e-81) (-4.7802e-81,-1.13699e-81) (-7.21054e-82,-3.69272e-81) (3.06471e-81,-6.77598e-82) (2.18342e-81,1.19186e-81) (-4.82607e-82,1.15561e-81) (-1.33643e-81,6.82023e-82) (-6.86855e-82,2.98568e-83) (-1.32541e-82,-4.59069e-82) (1.56682e-83,-4.68298e-82) (7.18375e-83,-2.3543e-82) (1.1568e-82,-6.74449e-83) (1.07479e-82,-9.16901e-84) (6.77189e-83,3.81211e-84) (3.3552e-83,6.44949e-84) (1.49741e-83,5.59401e-84) (6.58641e-84,3.3658e-84) (2.89031e-84,1.49617e-84) (1.22215e-84,4.84173e-85) (4.7466e-85,8.75002e-86) (1.59668e-85,-1.61675e-86) (4.30294e-86,-2.16551e-86) (8.04544e-87,-1.02644e-86) (5.04134e-88,-3.15164e-87) (-2.8063e-88,-6.51328e-88) (-1.23029e-88,-7.46531e-89) (-2.66355e-89,3.24164e-90) (-3.12046e-90,3.41903e-90) (2.4424e-92,7.4533e-91) 
  (1.05092e-94,6.54081e-94) (4.02029e-93,-3.08981e-93) (-3.39481e-92,-1.41353e-92) (3.5382e-92,2.51649e-91) (1.29086e-90,-1.06399e-90) (-9.97158e-90,-3.22041e-90) (1.7303e-89,5.98319e-89) (2.15341e-88,-2.7503e-88) (-1.83204e-87,-4.07701e-90) (5.72893e-87,6.78405e-87) (4.78075e-87,-3.89089e-86) (-1.21632e-85,9.6175e-86) (5.37716e-85,3.64347e-86) (-1.15957e-84,-1.11059e-84) (5.83359e-85,3.90784e-84) (3.45395e-84,-6.65108e-84) (-8.0551e-84,4.10572e-84) (-3.02547e-85,1.90037e-84) (2.88268e-83,8.96053e-84) (-5.32383e-83,-4.26658e-83) (6.36537e-83,3.76243e-83) (-1.31692e-82,5.92236e-83) (2.54131e-82,-1.61973e-82) (-1.72937e-82,2.26511e-82) (-2.20793e-82,-3.95834e-82) (5.33448e-82,4.54604e-82) (-5.26704e-82,1.42523e-82) (2.84061e-82,-9.41642e-82) (4.01909e-82,7.89283e-82) (-1.01742e-81,2.29128e-82) (2.91337e-82,-1.0119e-81) (9.61854e-82,6.39166e-82) (-6.50063e-82,6.8184e-82) (-6.58465e-82,-9.00019e-82) (6.59792e-82,-4.54881e-82) (5.16916e-82,6.50419e-82) (-4.77336e-82,4.2987e-82) (-4.87558e-82,-2.12919e-82) (1.46285e-82,-3.65939e-82) (3.28485e-82,-1.45065e-82) (1.06065e-82,1.19822e-82) (-4.11245e-83,1.95589e-82) (-5.92505e-83,9.20446e-83) (-5.843e-83,-1.4396e-83) (-4.81274e-83,-4.19728e-83) (-2.13904e-83,-3.0361e-83) (7.53844e-85,-1.89479e-83) (7.81069e-84,-1.22664e-83) (6.4215e-84,-6.97041e-84) (3.75476e-84,-3.15512e-84) (1.96386e-84,-1.19196e-84) (9.57778e-85,-4.3885e-85) (4.23489e-85,-1.86536e-85) (1.64012e-85,-9.1027e-86) (5.31896e-86,-4.4262e-86) (1.3085e-86,-1.9067e-86) (1.69235e-87,-6.77393e-87) (-3.5148e-88,-1.87077e-87) (-2.96198e-88,-3.64302e-88) (-9.94783e-89,-3.42552e-89) (-2.07011e-89,5.91965e-90) (-2.39653e-90,3.2618e-90) (4.83427e-92,7.01921e-91) (8.45757e-92,7.66844e-92) 
  (7.39313e-95,7.15841e-95) (2.10569e-94,-7.54806e-94) (-5.48248e-93,1.40628e-93) (2.76645e-92,2.74856e-92) (5.77609e-92,-2.49548e-91) (-1.50461e-90,5.47236e-91) (7.72865e-90,5.49943e-90) (-9.65746e-91,-5.28986e-89) (-2.11597e-88,1.7581e-88) (1.30011e-87,2.10735e-88) (-3.22806e-87,-4.72463e-87) (-3.71743e-87,2.1874e-86) (5.87135e-86,-4.71108e-86) (-2.17669e-85,-2.38117e-87) (4.06156e-85,3.16646e-85) (-2.59509e-85,-8.81065e-85) (-3.21964e-85,8.94591e-85) (-1.98391e-85,5.73788e-85) (4.03172e-84,-2.10047e-84) (-8.81089e-84,1.4158e-84) (8.36225e-84,-4.22167e-84) (-5.63938e-84,2.0536e-83) (6.47957e-84,-3.88143e-83) (1.1236e-83,3.30702e-83) (-6.36957e-83,-1.13428e-83) (8.70792e-83,-1.35183e-83) (-2.09876e-83,7.0264e-83) (-7.14773e-83,-1.10795e-82) (1.0954e-82,1.63062e-83) (-5.9342e-83,1.27986e-82) (-8.4465e-83,-1.08814e-82) (1.43377e-82,-4.90012e-83) (2.76243e-83,1.23919e-82) (-1.46597e-82,-4.50819e-84) (-3.1205e-84,-1.07512e-82) (1.11192e-82,-3.87241e-84) (1.18334e-83,8.32799e-83) (-6.38899e-83,3.82923e-83) (-2.89937e-83,-4.01609e-83) (1.23421e-83,-4.88585e-83) (2.12604e-83,-6.3042e-84) (1.67246e-83,1.97917e-83) (5.75665e-84,1.57775e-83) (-5.24394e-84,5.95637e-84) (-8.38251e-84,1.5702e-84) (-5.46497e-84,-3.17873e-85) (-2.23265e-84,-1.58849e-84) (-7.00788e-85,-1.82729e-84) (-1.87839e-85,-1.29717e-84) (-1.10024e-86,-6.97693e-85) (4.08474e-86,-3.26293e-85) (3.53721e-86,-1.45456e-85) (1.69556e-86,-6.33199e-86) (4.74324e-87,-2.62197e-86) (-4.65333e-90,-9.87616e-87) (-8.78442e-88,-3.1996e-87) (-5.82401e-88,-8.22381e-88) (-2.3822e-88,-1.40521e-88) (-6.86665e-89,-3.10018e-90) (-1.36098e-89,7.47752e-90) (-1.44235e-90,2.8619e-90) (1.11016e-91,5.97286e-91) (8.195e-92,6.7921e-92) (1.73605e-92,-1.16006e-93) 
  (1.57705e-95,2.05068e-96) (-4.35849e-95,-1.12388e-94) (-5.41913e-94,6.77639e-94) (5.91184e-93,7.88107e-94) (-1.6246e-92,-3.55656e-92) (-1.29006e-91,2.06905e-91) (1.43666e-90,-8.14609e-92) (-5.17112e-90,-6.06966e-90) (-7.22942e-90,4.04133e-89) (1.65031e-88,-1.01839e-88) (-8.03392e-88,-2.01249e-88) (1.69419e-87,2.64977e-87) (1.52845e-87,-1.02919e-86) (-2.14369e-86,1.97669e-86) (6.57827e-86,-6.65937e-87) (-9.55046e-86,-5.42887e-86) (3.52973e-86,8.44108e-86) (3.64525e-86,1.35959e-85) (1.94576e-85,-6.29346e-85) (-6.10343e-85,9.68395e-85) (1.04531e-85,-1.23139e-84) (1.71004e-84,2.54155e-84) (-3.15999e-84,-3.91432e-84) (4.28313e-84,1.02654e-84) (-6.97455e-84,5.76323e-84) (5.62308e-84,-9.28548e-84) (6.5944e-84,7.76563e-84) (-1.71791e-83,-2.33631e-84) (9.51013e-84,-1.02552e-83) (8.62267e-84,1.68346e-83) (-1.80387e-83,6.02152e-85) (6.23266e-84,-1.86854e-83) (1.60756e-83,6.39559e-84) (-1.20586e-83,1.46868e-83) (-1.24795e-83,-7.66331e-84) (8.3098e-84,-1.21549e-83) (1.00189e-83,4.73032e-84) (-9.0919e-85,1.02448e-83) (-6.30209e-84,5.75721e-85) (-4.21725e-84,-5.43985e-84) (6.0922e-85,-3.227e-84) (3.2756e-84,-2.10895e-85) (2.3637e-84,7.73279e-85) (4.09159e-85,1.03763e-84) (-5.01196e-85,1.0022e-84) (-5.28903e-85,5.85453e-85) (-3.7512e-85,1.39506e-85) (-2.55279e-85,-6.73581e-86) (-1.54792e-85,-9.10868e-86) (-7.72827e-86,-6.087e-86) (-3.27416e-86,-3.34955e-86) (-1.30739e-86,-1.67071e-86) (-5.48257e-87,-7.45474e-87) (-2.44954e-87,-2.86374e-87) (-1.08032e-87,-8.95448e-88) (-4.3034e-88,-1.98696e-88) (-1.44211e-88,-1.33674e-89) (-3.79729e-89,1.26137e-89) (-6.98058e-90,7.18309e-90) (-5.25542e-91,2.21915e-90) (1.6729e-91,4.44084e-91) (7.64603e-92,4.8814e-92) (1.59096e-92,-1.90488e-93) (1.69958e-93,-2.01992e-93) 
  (2.13442e-96,-1.19059e-96) (-1.56392e-95,-9.79658e-96) (-3.84645e-96,1.32434e-94) (7.89523e-94,-4.5071e-94) (-5.26807e-93,-2.76608e-93) (4.09492e-93,3.67788e-92) (1.61035e-91,-1.45994e-91) (-1.1775e-90,-2.05445e-91) (3.06888e-90,5.25623e-90) (8.36476e-90,-2.7071e-89) (-1.05152e-88,5.53674e-89) (4.26578e-88,1.13964e-88) (-8.06846e-88,-1.17187e-87) (-2.58811e-88,3.8488e-87) (5.40601e-87,-6.3654e-87) (-1.23563e-86,3.1907e-87) (6.64981e-87,3.39511e-87) (2.17457e-86,1.4686e-86) (-4.42598e-86,-8.12486e-86) (4.3222e-86,1.37849e-85) (-1.36005e-85,-1.02423e-85) (4.26293e-85,5.61635e-86) (-6.30057e-85,-2.33136e-86) (4.10987e-85,-4.0794e-85) (-3.22576e-86,1.23773e-84) (-4.45775e-85,-1.23547e-84) (1.43272e-84,-1.36041e-85) (-1.6689e-84,1.48832e-84) (-4.20166e-85,-1.74929e-84) (2.46162e-84,4.85288e-85) (-1.32194e-84,1.9686e-84) (-1.44172e-84,-2.09019e-84) (1.98098e-84,-1.30387e-84) (5.69001e-85,2.36043e-84) (-1.83025e-84,8.37417e-85) (-6.46829e-85,-1.81468e-84) (1.25263e-84,-7.72788e-85) (1.0501e-84,9.23051e-85) (-3.42809e-85,7.59819e-85) (-9.16604e-85,1.17517e-87) (-3.74857e-85,-3.28861e-85) (2.10335e-85,-3.5099e-85) (2.97904e-85,-1.95995e-85) (1.63556e-85,2.10982e-86) (6.74875e-86,1.29115e-85) (1.76862e-86,1.0995e-85) (-1.49987e-86,5.65764e-86) (-2.74293e-86,2.30634e-86) (-2.2758e-86,8.85608e-87) (-1.34061e-86,3.02606e-87) (-6.60047e-87,6.61777e-88) (-2.99756e-87,-1.42985e-89) (-1.30113e-87,-5.16626e-89) (-5.30608e-88,1.31926e-89) (-1.94989e-88,3.69508e-89) (-6.1028e-89,2.86315e-89) (-1.48684e-89,1.44387e-89) (-2.21874e-90,5.32021e-90) (1.09488e-91,1.44901e-90) (1.89649e-91,2.74112e-91) (6.48796e-92,2.60315e-92) (1.30471e-92,-3.36232e-93) (1.4315e-93,-1.926e-93) (-4.22532e-95,-3.96379e-94) 
  (1.53862e-97,-3.40231e-97) (-2.80225e-96,2.30242e-97) (1.1678e-95,1.64258e-95) (5.35536e-95,-1.27334e-94) (-8.88215e-94,1.60784e-94) (3.951e-93,3.96314e-93) (4.86816e-93,-3.2319e-92) (-1.54173e-91,8.926e-92) (8.47194e-91,2.92055e-91) (-1.68583e-90,-3.74492e-90) (-5.82747e-90,1.58636e-89) (5.43481e-89,-2.85252e-89) (-1.88015e-88,-4.09069e-89) (3.22389e-88,3.86978e-88) (-6.69977e-89,-1.03393e-87) (-7.42332e-88,1.22123e-87) (3.9511e-88,-3.0337e-90) (4.32346e-87,-6.89912e-88) (-1.22141e-86,-3.32039e-87) (1.67324e-86,6.69321e-87) (-2.28215e-86,7.95911e-87) (4.4761e-86,-3.83876e-86) (-5.2288e-86,5.73736e-86) (-1.66811e-86,-7.74283e-86) (1.21265e-85,1.13058e-85) (-1.49498e-85,-4.75949e-86) (1.05914e-85,-1.73739e-85) (7.29238e-87,2.82921e-85) (-2.22387e-85,-8.10545e-86) (2.50225e-85,-2.13578e-85) (1.08517e-85,2.92981e-85) (-3.24933e-85,-1.05635e-86) (1.33721e-86,-3.24792e-85) (2.82936e-85,1.18281e-85) (-4.85281e-86,2.73059e-85) (-2.40109e-85,-6.83039e-86) (4.72524e-87,-1.97171e-85) (1.82645e-85,-4.04297e-86) (6.71625e-86,9.17762e-86) (-7.17318e-86,9.53043e-86) (-7.25511e-86,1.98584e-86) (-2.29139e-86,-4.54055e-86) (4.4803e-87,-4.94695e-86) (1.56119e-86,-1.93897e-86) (1.87672e-86,2.2235e-87) (1.34339e-86,7.57383e-87) (5.35096e-87,6.61592e-87) (4.48934e-88,4.8858e-87) (-9.37835e-88,3.16439e-87) (-8.40209e-88,1.70745e-87) (-5.08029e-88,7.83103e-88) (-2.63571e-88,3.297e-88) (-1.19431e-88,1.38217e-88) (-4.54467e-89,5.89914e-89) (-1.34667e-89,2.44865e-89) (-2.45198e-90,9.22288e-90) (1.89002e-91,2.94666e-90) (3.67815e-91,7.40571e-91) (1.67455e-91,1.26605e-91) (4.81167e-92,6.08901e-93) (9.22991e-93,-4.45231e-93) (9.47843e-94,-1.75039e-93) (-6.21399e-95,-3.52005e-94) (-4.73872e-95,-3.66183e-95) 
  (-1.20062e-98,-5.5431e-98) (-3.19097e-97,2.8296e-97) (2.91647e-96,9.11118e-97) (-5.37284e-96,-2.02282e-95) (-9.04942e-95,1.02219e-94) (8.38076e-94,9.16845e-95) (-2.51644e-93,-4.19338e-93) (-8.88572e-93,2.48488e-92) (1.21487e-91,-4.89585e-92) (-5.38855e-91,-2.41192e-91) (8.96296e-91,2.20634e-90) (2.81381e-90,-7.96416e-90) (-2.20327e-89,1.32829e-89) (6.44619e-89,7.20857e-90) (-9.35533e-89,-8.43997e-89) (3.45128e-89,1.48414e-88) (1.32809e-89,3.94678e-89) (4.08875e-88,-5.46168e-88) (-1.44337e-87,8.83955e-88) (1.93135e-87,-1.12798e-87) (-9.91965e-88,3.32408e-87) (2.04703e-88,-7.90897e-87) (1.39273e-87,9.31732e-87) (-1.02681e-86,-4.20869e-87) (2.1637e-86,-2.00752e-87) (-1.49814e-86,1.11604e-86) (-9.87788e-87,-2.67214e-86) (2.76336e-86,2.1774e-86) (-2.57364e-86,1.8647e-86) (-1.64232e-87,-4.26002e-86) (3.97324e-86,1.10766e-86) (-2.53505e-86,3.27931e-86) (-3.45563e-86,-2.77459e-86) (3.25619e-86,-2.04471e-86) (2.66703e-86,2.7158e-86) (-2.48605e-86,2.03565e-86) (-2.1876e-86,-1.51275e-86) (9.80409e-87,-2.26281e-86) (1.58612e-86,-1.56793e-87) (4.45343e-87,1.45573e-86) (-3.81049e-87,1.04318e-86) (-6.4213e-87,-3.52285e-88) (-4.90347e-87,-4.62781e-87) (-1.11518e-87,-3.57453e-87) (1.57832e-87,-1.90135e-87) (1.94088e-87,-8.01254e-88) (1.22328e-87,-4.41123e-89) (5.89929e-88,3.33703e-88) (2.62536e-88,3.5839e-88) (1.10707e-88,2.36669e-88) (4.09379e-89,1.23863e-88) (1.32535e-89,5.76993e-89) (4.71805e-90,2.5105e-89) (2.41762e-90,1.01249e-89) (1.45086e-90,3.64001e-90) (7.74514e-91,1.09952e-90) (3.35464e-91,2.50603e-91) (1.14338e-91,2.95327e-92) (2.95869e-92,-6.0549e-93) (5.30417e-93,-4.60984e-93) (4.2507e-94,-1.43368e-93) (-9.43027e-95,-2.76972e-94) (-4.42805e-95,-2.90325e-95) (-8.84695e-96,1.33734e-96) 
  (-6.46118e-99,-5.62819e-99) (-1.26901e-98,6.31882e-98) (4.33742e-97,-1.59034e-97) (-2.52075e-96,-1.91109e-96) (-1.0793e-96,2.05587e-95) (1.06216e-94,-6.87205e-95) (-6.87463e-94,-2.39402e-94) (1.38317e-93,3.62932e-93) (8.57169e-93,-1.69567e-92) (-8.0129e-92,2.5694e-92) (3.00337e-91,1.42565e-91) (-4.60409e-91,-1.05434e-90) (-9.0092e-91,3.27835e-90) (6.51952e-90,-5.02711e-90) (-1.49641e-89,6.29307e-91) (1.2773e-89,8.07707e-90) (9.57294e-90,1.13755e-89) (-1.39796e-89,-1.00415e-88) (-4.34448e-89,2.17598e-88) (3.06232e-89,-2.76938e-88) (2.89282e-88,4.02933e-88) (-7.52825e-88,-7.17574e-88) (9.88638e-88,5.55004e-88) (-1.3376e-87,8.11964e-88) (1.65526e-87,-2.24561e-87) (1.18543e-88,2.24942e-87) (-3.70903e-87,-1.29274e-87) (4.19652e-87,-9.59424e-88) (6.91744e-89,4.32349e-87) (-4.43255e-87,-3.19645e-87) (4.27396e-87,-3.37988e-87) (1.55542e-87,5.04816e-87) (-5.8011e-87,1.47712e-87) (1.55571e-88,-4.81634e-87) (5.12264e-87,-7.56957e-88) (3.80269e-88,4.10968e-87) (-3.34276e-87,1.3267e-87) (-1.66284e-87,-2.74711e-87) (1.00546e-87,-2.02524e-87) (1.82667e-87,5.8118e-88) (8.79743e-88,1.33386e-87) (-4.41235e-88,7.21095e-88) (-8.8369e-88,1.41911e-88) (-5.26538e-88,-1.73063e-88) (-1.03811e-88,-3.12217e-88) (7.37301e-89,-2.7206e-88) (1.00506e-88,-1.4188e-88) (8.50926e-89,-4.07032e-89) (5.96961e-89,5.81035e-91) (3.46313e-89,8.26135e-90) (1.69637e-89,6.32354e-90) (7.45936e-90,3.56421e-90) (3.14791e-90,1.6644e-90) (1.30925e-90,6.23487e-91) (5.21577e-91,1.65915e-91) (1.88094e-91,1.54779e-92) (5.7622e-92,-1.31806e-92) (1.38043e-92,-9.55327e-93) (2.14429e-93,-3.75685e-93) (1.27223e-95,-1.014e-93) (-1.13002e-94,-1.85608e-94) (-3.91598e-95,-1.72877e-95) (-7.58198e-96,1.83762e-96) (-7.62483e-97,1.08858e-96) 
  (-1.27194e-99,-8.31694e-101) (4.26482e-99,8.60884e-99) (3.62676e-98,-5.86707e-98) (-4.72091e-97,1.21365e-98) (1.8111e-96,2.47332e-96) (5.54795e-96,-1.7893e-95) (-9.95116e-95,3.89418e-95) (4.98193e-94,2.6319e-94) (-7.1112e-94,-2.6211e-93) (-5.82899e-93,1.02792e-92) (4.35114e-92,-1.40473e-92) (-1.42529e-91,-5.91984e-92) (2.14469e-91,3.86605e-91) (1.33155e-91,-1.01662e-90) (-1.15987e-90,1.28208e-90) (1.28713e-90,-3.08051e-91) (3.11944e-90,5.00637e-91) (-1.1713e-89,-8.53786e-90) (1.73087e-89,2.27004e-89) (-2.6511e-89,-2.30726e-89) (6.9889e-89,3.29572e-90) (-1.33466e-88,1.2126e-89) (1.23489e-88,-5.83086e-89) (-2.32051e-89,2.17926e-88) (-7.92192e-89,-3.42026e-88) (2.47212e-88,1.32484e-88) (-4.54086e-88,2.77302e-88) (2.10971e-88,-4.76218e-88) (4.88845e-88,3.32772e-88) (-6.61998e-88,2.10274e-88) (-3.80097e-89,-7.18418e-88) (6.48842e-88,1.90914e-88) (-2.99822e-88,7.41031e-88) (-5.07409e-88,-3.37403e-88) (3.16945e-88,-6.19678e-88) (4.74116e-88,2.41121e-88) (-9.63834e-89,4.75835e-88) (-4.13847e-88,-1.8011e-89) (-1.65446e-88,-2.74051e-88) (1.82987e-88,-1.55359e-88) (2.23445e-88,1.05342e-89) (6.04165e-89,9.94869e-89) (-5.20152e-89,1.04195e-88) (-6.47559e-89,4.73523e-89) (-4.37696e-89,-9.4687e-90) (-2.34359e-89,-2.9089e-89) (-7.49016e-90,-2.31376e-89) (2.03188e-90,-1.30015e-89) (4.71554e-90,-6.47262e-90) (3.72652e-90,-3.03756e-90) (2.11873e-90,-1.3051e-90) (1.02389e-90,-5.14258e-91) (4.49462e-91,-2.03109e-91) (1.79816e-91,-8.90626e-92) (6.31619e-92,-4.20694e-92) (1.82184e-92,-1.89279e-92) (3.73447e-93,-7.37898e-93) (2.29623e-94,-2.35238e-93) (-2.04934e-94,-5.78185e-94) (-1.07735e-94,-9.68458e-95) (-3.07443e-95,-5.61496e-96) (-5.65728e-96,2.52185e-96) (-5.5132e-97,9.92653e-97) (3.98043e-98,1.90656e-97) ]
